module wallypipelinedcorewrapper (
	clk,
	reset,
	MTimerInt,
	MExtInt,
	SExtInt,
	MSwInt,
	MTIME_CLINT,
	HRDATA,
	HREADY,
	HRESP,
	HCLK,
	HRESETn,
	HADDR,
	HWDATA,
	HWSTRB,
	HWRITE,
	HSIZE,
	HBURST,
	HPROT,
	HTRANS,
	HMASTLOCK,
	ExternalStall
);
	input wire clk;
	input wire reset;
	input wire MTimerInt;
	input wire MExtInt;
	input wire SExtInt;
	input wire MSwInt;
	input wire [63:0] MTIME_CLINT;
	localparam XLEN = 32'd64;
	localparam AHBW = XLEN;
	localparam ASID_BASE = 32'd44;
	localparam ASID_BITS = 32'd16;
	localparam [0:0] ZAAMO_SUPPORTED = 1;
	localparam [0:0] ZALRSC_SUPPORTED = 1;
	localparam [0:0] A_SUPPORTED = ZAAMO_SUPPORTED & ZALRSC_SUPPORTED;
	localparam D_BIAS = 32'd1023;
	localparam [0:0] D_SUPPORTED = 1;
	localparam Q_BIAS = 32'd16383;
	localparam [0:0] Q_SUPPORTED = 0;
	localparam S_BIAS = 32'd127;
	localparam BIAS = (Q_SUPPORTED ? Q_BIAS : (D_SUPPORTED ? D_BIAS : S_BIAS));
	localparam D_LEN = 32'd64;
	localparam Q_LEN = 32'd128;
	localparam S_LEN = 32'd32;
	localparam FLEN = (Q_SUPPORTED ? Q_LEN : (D_SUPPORTED ? D_LEN : S_LEN));
	localparam H_BIAS = 32'd15;
	localparam BIAS1 = (FLEN > D_LEN ? D_BIAS : (FLEN > S_LEN ? S_BIAS : H_BIAS));
	localparam H_LEN = 32'd16;
	localparam LEN1 = (FLEN > D_LEN ? D_LEN : (FLEN > S_LEN ? S_LEN : H_LEN));
	localparam BIAS2 = (LEN1 > S_LEN ? S_BIAS : H_BIAS);
	localparam [0:0] BIGENDIAN_SUPPORTED = 1;
	localparam [63:0] BOOTROM_BASE = 64'h0000000000001000;
	localparam [0:0] BOOTROM_PRELOAD = 1'b0;
	localparam [63:0] BOOTROM_RANGE = 64'h0000000000000fff;
	localparam [0:0] BOOTROM_SUPPORTED = 1;
	localparam BPRED_NUM_LHR = 32'd6;
	localparam BPRED_SIZE = 32'd10;
	localparam [0:0] BPRED_SUPPORTED = 1;
	localparam BPRED_TYPE = 32'd1;
	localparam BTB_SIZE = 32'd10;
	localparam [0:0] BURST_EN = 1;
	localparam [0:0] BUS_SUPPORTED = 1;
	localparam [0:0] ZBA_SUPPORTED = 1;
	localparam [0:0] ZBB_SUPPORTED = 1;
	localparam [0:0] ZBS_SUPPORTED = 1;
	localparam [0:0] B_SUPPORTED = (ZBA_SUPPORTED & ZBB_SUPPORTED) & ZBS_SUPPORTED;
	localparam CACHE_SRAMLEN = 32'd128;
	localparam [63:0] CLINT_BASE = 64'h0000000002000000;
	localparam [63:0] CLINT_RANGE = 64'h000000000000ffff;
	localparam [0:0] CLINT_SUPPORTED = 1;
	localparam COUNTERS = 12'd32;
	localparam D_NF = 32'd52;
	localparam Q_NF = 32'd112;
	localparam S_NF = 32'd23;
	localparam NF = (Q_SUPPORTED ? Q_NF : (D_SUPPORTED ? D_NF : S_NF));
	localparam BASECVTLEN = (XLEN > NF ? XLEN : NF);
	localparam [0:0] ZFA_SUPPORTED = 1;
	localparam CVTLEN = (ZFA_SUPPORTED & D_SUPPORTED ? (BASECVTLEN > 32'd84 ? BASECVTLEN : 32'd84) : BASECVTLEN);
	localparam [0:0] F_SUPPORTED = 1;
	localparam [0:0] ZCA_SUPPORTED = 1;
	localparam [0:0] ZCD_SUPPORTED = 1;
	localparam [0:0] ZCF_SUPPORTED = 0;
	localparam [0:0] C_SUPPORTED = (ZCA_SUPPORTED & (D_SUPPORTED ? ZCD_SUPPORTED : 1)) & (F_SUPPORTED ? 1 : 1);
	localparam DCACHE_LINELENINBITS = 32'd512;
	localparam DCACHE_NUMWAYS = 32'd4;
	localparam [0:0] DCACHE_SUPPORTED = 1;
	localparam DCACHE_WAYSIZEINBYTES = 32'd4096;
	localparam FPDIVMINb = NF + 2;
	localparam [0:0] IDIV_ON_FPU = 1;
	localparam DIVMINb = ((FPDIVMINb < XLEN) & IDIV_ON_FPU ? XLEN : FPDIVMINb);
	localparam RADIX = 32'd4;
	localparam LOGR = 2;
	localparam RESBITS = DIVMINb + LOGR;
	localparam DIVCOPIES = 32'd4;
	localparam RK = 8;
	localparam FPDUR = ((RESBITS - 1) / RK) + 1;
	localparam DIVb = (FPDUR * RK) - LOGR;
	localparam DIVBLEN = $clog2(DIVb + 1);
	localparam [63:0] DTIM_BASE = 64'h0000000080000000;
	localparam [63:0] DTIM_RANGE = 64'h00000000007fffff;
	localparam [0:0] DTIM_SUPPORTED = 0;
	localparam DTLB_ENTRIES = 32'd32;
	localparam DURLEN = $clog2(FPDUR);
	localparam D_FMT = 2'd1;
	localparam D_NE = 32'd11;
	localparam [63:0] EXT_MEM_BASE = 64'h0000000080000000;
	localparam [63:0] EXT_MEM_RANGE = 64'h0000000007ffffff;
	localparam [0:0] EXT_MEM_SUPPORTED = 0;
	localparam [0:0] E_SUPPORTED = 0;
	localparam FMALEN = (3 * NF) + 6;
	localparam FMT = (Q_SUPPORTED ? 2'd3 : (D_SUPPORTED ? 2'd1 : 2'd0));
	localparam FMT1 = (FLEN > D_LEN ? 2'd1 : (FLEN > S_LEN ? 2'd0 : 2'd2));
	localparam FMT2 = (LEN1 > S_LEN ? 2'd0 : 2'd2);
	localparam [0:0] ZFH_SUPPORTED = 1;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	localparam FPSIZES = ((sv2v_cast_32(Q_SUPPORTED) + sv2v_cast_32(D_SUPPORTED)) + sv2v_cast_32(F_SUPPORTED)) + sv2v_cast_32(ZFH_SUPPORTED);
	localparam FMTBITS = sv2v_cast_32(FPSIZES >= 3) + 1;
	localparam [63:0] GPIO_BASE = 64'h0000000010060000;
	localparam [0:0] GPIO_LOOPBACK_TEST = 1;
	localparam [63:0] GPIO_RANGE = 64'h00000000000000ff;
	localparam [0:0] GPIO_SUPPORTED = 1;
	localparam H_FMT = 2'd2;
	localparam H_NE = 32'd5;
	localparam H_NF = 32'd10;
	localparam ICACHE_LINELENINBITS = 32'd512;
	localparam ICACHE_NUMWAYS = 32'd4;
	localparam [0:0] ICACHE_SUPPORTED = 1;
	localparam ICACHE_WAYSIZEINBYTES = 32'd4096;
	localparam IDIV_BITSPERCYCLE = 32'd4;
	localparam [0:0] IEEE754 = 0;
	localparam INSTR_CLASS_PRED = 1;
	localparam INTRESBITS = 66;
	localparam INTFPDUR = 9;
	localparam INTDIVb = 70;
	localparam [63:0] IROM_BASE = 64'h0000000080000000;
	localparam [63:0] IROM_RANGE = 64'h00000000007fffff;
	localparam [0:0] IROM_SUPPORTED = 0;
	localparam ITLB_ENTRIES = 32'd32;
	localparam [0:0] I_SUPPORTED = !E_SUPPORTED;
	localparam LEN2 = (LEN1 > S_LEN ? S_LEN : H_LEN);
	localparam LLEN = ($unsigned(FLEN) > $unsigned(XLEN) ? $unsigned(FLEN) : $unsigned(XLEN));
	localparam LOGCVTLEN = $unsigned($clog2(CVTLEN + 1));
	localparam LOGFLEN = $clog2(FLEN);
	localparam NORMSHIFTSZ = ((((CVTLEN + NF) + 1) > (((DIVb + 1) + NF) + 1) ? (CVTLEN + NF) + 1 : ((DIVb + 1) + NF) + 1) > (FMALEN + 2) ? (((CVTLEN + NF) + 1) > (((DIVb + 1) + NF) + 1) ? (CVTLEN + NF) + 1 : ((DIVb + 1) + NF) + 1) : FMALEN + 2);
	localparam LOGNORMSHIFTSZ = $clog2(NORMSHIFTSZ);
	localparam LOG_XLEN = 32'd6;
	localparam [0:0] M_SUPPORTED = 1;
	localparam [0:0] S_SUPPORTED = 1;
	localparam [0:0] U_SUPPORTED = 1;
	localparam MISA = {11'b00000000000, U_SUPPORTED, 1'b0, S_SUPPORTED, 1'b0, Q_SUPPORTED, 3'b000, M_SUPPORTED, 3'b000, I_SUPPORTED, 2'b00, F_SUPPORTED, E_SUPPORTED, D_SUPPORTED, C_SUPPORTED, B_SUPPORTED, A_SUPPORTED};
	localparam M_MODE = 2'b11;
	localparam Q_NE = 32'd15;
	localparam S_NE = 32'd8;
	localparam NE = (Q_SUPPORTED ? Q_NE : (D_SUPPORTED ? D_NE : S_NE));
	localparam NE1 = (FLEN > D_LEN ? D_NE : (FLEN > S_LEN ? S_NE : H_NE));
	localparam NE2 = (LEN1 > S_LEN ? S_NE : H_NE);
	localparam NF1 = (FLEN > D_LEN ? D_NF : (FLEN > S_LEN ? S_NF : H_NF));
	localparam NF2 = (LEN1 > S_LEN ? S_NF : H_NF);
	localparam NO_TRANSLATE = 4'd0;
	localparam PA_BITS = 32'd56;
	localparam [63:0] PLIC_BASE = 64'h000000000c000000;
	localparam PLIC_GPIO_ID = 32'd3;
	localparam PLIC_NUM_SRC = 32'd10;
	localparam PLIC_NUM_SRC_LT_32 = 1'd1;
	localparam [63:0] PLIC_RANGE = 64'h0000000003ffffff;
	localparam PLIC_SDC_ID = 32'd9;
	localparam PLIC_SPI_ID = 32'd6;
	localparam [0:0] PLIC_SUPPORTED = 1;
	localparam PLIC_UART_ID = 32'd10;
	localparam PMP_ENTRIES = 32'd16;
	localparam PMPCFG_ENTRIES = PMP_ENTRIES / 32'd8;
	localparam PPN_BITS = 32'd44;
	localparam Q_FMT = 2'd3;
	localparam RAM_LATENCY = 32'b00000000000000000000000000000000;
	localparam RAS_SIZE = 32'd16;
	localparam [63:0] RESET_VECTOR = 64'h0000000080000000;
	localparam [63:0] SDC_BASE = 64'h0000000000013000;
	localparam [63:0] SDC_RANGE = 64'h0000000000000fff;
	localparam [0:0] SDC_SUPPORTED = 0;
	localparam [63:0] SPI_BASE = 64'h0000000010040000;
	localparam [0:0] SPI_LOOPBACK_TEST = 1;
	localparam [63:0] SPI_RANGE = 64'h0000000000000fff;
	localparam [0:0] SPI_SUPPORTED = 1;
	localparam [0:0] SSTC_SUPPORTED = 1;
	localparam SV32 = 4'd1;
	localparam SV39 = 4'd8;
	localparam SV48 = 4'd9;
	localparam [0:0] SVADU_SUPPORTED = 1;
	localparam [0:0] SVINVAL_SUPPORTED = 1;
	localparam SVMODE_BITS = 32'd4;
	localparam [0:0] SVNAPOT_SUPPORTED = 1;
	localparam [0:0] SVPBMT_SUPPORTED = 1;
	localparam S_FMT = 2'd0;
	localparam S_MODE = 2'b01;
	localparam [63:0] UART_BASE = 64'h0000000010000000;
	localparam UART_PRESCALE = 32'd1;
	localparam [63:0] UART_RANGE = 64'h0000000000000007;
	localparam [0:0] UART_SUPPORTED = 1;
	localparam [63:0] UNCORE_RAM_BASE = 64'h0000000080000000;
	localparam [0:0] UNCORE_RAM_PRELOAD = 1'b0;
	localparam [63:0] UNCORE_RAM_RANGE = 64'h0000000007ffffff;
	localparam [0:0] UNCORE_RAM_SUPPORTED = 1;
	localparam [0:0] USE_SRAM = 0;
	localparam U_MODE = 2'b00;
	localparam [0:0] VECTORED_INTERRUPTS_SUPPORTED = 1;
	localparam [0:0] VIRTMEM_SUPPORTED = 1;
	localparam VPN_SEGMENT_BITS = 32'd9;
	localparam VPN_BITS = 36;
	localparam WFI_TIMEOUT_BIT = 32'd16;
	localparam [0:0] ZBC_SUPPORTED = 1;
	localparam [0:0] ZBKB_SUPPORTED = 1;
	localparam [0:0] ZBKC_SUPPORTED = 1;
	localparam [0:0] ZBKX_SUPPORTED = 1;
	localparam [0:0] ZCB_SUPPORTED = 1;
	localparam [0:0] ZICBOM_SUPPORTED = 1;
	localparam [0:0] ZICBOP_SUPPORTED = 1;
	localparam [0:0] ZICBOZ_SUPPORTED = 1;
	localparam [0:0] ZICCLSM_SUPPORTED = 1;
	localparam [0:0] ZICNTR_SUPPORTED = 1;
	localparam [0:0] ZICOND_SUPPORTED = 1;
	localparam [0:0] ZICSR_SUPPORTED = 1;
	localparam [0:0] ZIFENCEI_SUPPORTED = 1;
	localparam [0:0] ZIHPM_SUPPORTED = 1;
	localparam [0:0] ZKND_SUPPORTED = 1;
	localparam [0:0] ZKNE_SUPPORTED = 1;
	localparam [0:0] ZKNH_SUPPORTED = 1;
	localparam [0:0] ZKN_SUPPORTED = ((((ZBKB_SUPPORTED & ZBKC_SUPPORTED) & ZBKX_SUPPORTED) & ZKND_SUPPORTED) & ZKNE_SUPPORTED) & ZKNH_SUPPORTED;
	localparam [0:0] ZMMUL_SUPPORTED = 1;
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	localparam [4216:0] P = {sv2v_cast_32_signed(XLEN), IEEE754, sv2v_cast_32_signed(MISA), sv2v_cast_32_signed(AHBW), sv2v_cast_32_signed(RAM_LATENCY), BURST_EN, ZICSR_SUPPORTED, ZIFENCEI_SUPPORTED, COUNTERS, ZICNTR_SUPPORTED, ZIHPM_SUPPORTED, ZFH_SUPPORTED, ZFA_SUPPORTED, SSTC_SUPPORTED, VIRTMEM_SUPPORTED, VECTORED_INTERRUPTS_SUPPORTED, BIGENDIAN_SUPPORTED, SVADU_SUPPORTED, ZMMUL_SUPPORTED, ZICBOM_SUPPORTED, ZICBOZ_SUPPORTED, ZICBOP_SUPPORTED, ZICCLSM_SUPPORTED, ZICOND_SUPPORTED, SVPBMT_SUPPORTED, SVNAPOT_SUPPORTED, SVINVAL_SUPPORTED, ZAAMO_SUPPORTED, ZALRSC_SUPPORTED, BUS_SUPPORTED, DCACHE_SUPPORTED, ICACHE_SUPPORTED, sv2v_cast_32_signed(ITLB_ENTRIES), sv2v_cast_32_signed(DTLB_ENTRIES), sv2v_cast_32_signed(DCACHE_NUMWAYS), sv2v_cast_32_signed(DCACHE_WAYSIZEINBYTES), sv2v_cast_32_signed(DCACHE_LINELENINBITS), sv2v_cast_32_signed(ICACHE_NUMWAYS), sv2v_cast_32_signed(ICACHE_WAYSIZEINBYTES), sv2v_cast_32_signed(ICACHE_LINELENINBITS), sv2v_cast_32_signed(CACHE_SRAMLEN), sv2v_cast_32_signed(IDIV_BITSPERCYCLE), IDIV_ON_FPU, sv2v_cast_32_signed(PMP_ENTRIES), RESET_VECTOR, sv2v_cast_32_signed(WFI_TIMEOUT_BIT), DTIM_SUPPORTED, DTIM_BASE, DTIM_RANGE, IROM_SUPPORTED, IROM_BASE, IROM_RANGE, BOOTROM_SUPPORTED, BOOTROM_BASE, BOOTROM_RANGE, BOOTROM_PRELOAD, UNCORE_RAM_SUPPORTED, UNCORE_RAM_BASE, UNCORE_RAM_RANGE, UNCORE_RAM_PRELOAD, EXT_MEM_SUPPORTED, EXT_MEM_BASE, EXT_MEM_RANGE, CLINT_SUPPORTED, CLINT_BASE, CLINT_RANGE, GPIO_SUPPORTED, GPIO_BASE, GPIO_RANGE, UART_SUPPORTED, UART_BASE, UART_RANGE, PLIC_SUPPORTED, PLIC_BASE, PLIC_RANGE, SDC_SUPPORTED, SDC_BASE, SDC_RANGE, SPI_SUPPORTED, SPI_BASE, SPI_RANGE, GPIO_LOOPBACK_TEST, SPI_LOOPBACK_TEST, sv2v_cast_32_signed(UART_PRESCALE), sv2v_cast_32_signed(PLIC_NUM_SRC), PLIC_NUM_SRC_LT_32, sv2v_cast_32_signed(PLIC_GPIO_ID), sv2v_cast_32_signed(PLIC_UART_ID), sv2v_cast_32_signed(PLIC_SPI_ID), sv2v_cast_32_signed(PLIC_SDC_ID), BPRED_SUPPORTED, BPRED_TYPE, sv2v_cast_32_signed(BPRED_NUM_LHR), sv2v_cast_32_signed(BPRED_SIZE), sv2v_cast_32_signed(BTB_SIZE), sv2v_cast_32_signed(RAS_SIZE), sv2v_cast_1(INSTR_CLASS_PRED), sv2v_cast_32_signed(RADIX), sv2v_cast_32_signed(DIVCOPIES), ZBA_SUPPORTED, ZBB_SUPPORTED, ZBC_SUPPORTED, ZBS_SUPPORTED, ZCA_SUPPORTED, ZCB_SUPPORTED, ZCD_SUPPORTED, ZCF_SUPPORTED, ZBKB_SUPPORTED, ZBKC_SUPPORTED, ZBKX_SUPPORTED, ZKND_SUPPORTED, ZKNE_SUPPORTED, ZKNH_SUPPORTED, ZKN_SUPPORTED, USE_SRAM, M_MODE, S_MODE, U_MODE, sv2v_cast_32_signed(VPN_SEGMENT_BITS), VPN_BITS, sv2v_cast_32_signed(PPN_BITS), sv2v_cast_32_signed(PA_BITS), sv2v_cast_32_signed(SVMODE_BITS), sv2v_cast_32_signed(ASID_BASE), sv2v_cast_32_signed(ASID_BITS), NO_TRANSLATE, SV32, SV39, SV48, A_SUPPORTED, B_SUPPORTED, C_SUPPORTED, D_SUPPORTED, E_SUPPORTED, F_SUPPORTED, I_SUPPORTED, M_SUPPORTED, Q_SUPPORTED, S_SUPPORTED, U_SUPPORTED, sv2v_cast_32_signed(LOG_XLEN), sv2v_cast_32_signed(PMPCFG_ENTRIES), sv2v_cast_32_signed(Q_LEN), sv2v_cast_32_signed(Q_NE), sv2v_cast_32_signed(Q_NF), sv2v_cast_32_signed(Q_BIAS), Q_FMT, sv2v_cast_32_signed(D_LEN), sv2v_cast_32_signed(D_NE), sv2v_cast_32_signed(D_NF), sv2v_cast_32_signed(D_BIAS), D_FMT, sv2v_cast_32_signed(S_LEN), sv2v_cast_32_signed(S_NE), sv2v_cast_32_signed(S_NF), sv2v_cast_32_signed(S_BIAS), S_FMT, sv2v_cast_32_signed(H_LEN), sv2v_cast_32_signed(H_NE), sv2v_cast_32_signed(H_NF), sv2v_cast_32_signed(H_BIAS), H_FMT, sv2v_cast_32_signed(FLEN), LOGFLEN, sv2v_cast_32_signed(NE), sv2v_cast_32_signed(NF), FMT, sv2v_cast_32_signed(BIAS), sv2v_cast_32_signed(FPSIZES), sv2v_cast_32_signed(FMTBITS), sv2v_cast_32_signed(LEN1), sv2v_cast_32_signed(NE1), sv2v_cast_32_signed(NF1), FMT1, sv2v_cast_32_signed(BIAS1), sv2v_cast_32_signed(LEN2), sv2v_cast_32_signed(NE2), sv2v_cast_32_signed(NF2), FMT2, sv2v_cast_32_signed(BIAS2), sv2v_cast_32_signed(CVTLEN), sv2v_cast_32_signed(LLEN), sv2v_cast_32_signed(LOGCVTLEN), sv2v_cast_32_signed(NORMSHIFTSZ), LOGNORMSHIFTSZ, sv2v_cast_32_signed(FMALEN), LOGR, RK, sv2v_cast_32_signed(FPDUR), DURLEN, sv2v_cast_32_signed(DIVb), DIVBLEN, INTDIVb};
	input wire [$signed(P[4151-:32]) - 1:0] HRDATA;
	input wire HREADY;
	input wire HRESP;
	output wire HCLK;
	output wire HRESETn;
	output wire [$signed(P[1640-:32]) - 1:0] HADDR;
	output wire [$signed(P[4151-:32]) - 1:0] HWDATA;
	output wire [($signed(P[4216-:32]) / 8) - 1:0] HWSTRB;
	output wire HWRITE;
	output wire [2:0] HSIZE;
	output wire [2:0] HBURST;
	output wire [3:0] HPROT;
	output wire [1:0] HTRANS;
	output wire HMASTLOCK;
	input wire ExternalStall;
	wallypipelinedcore #(.P(P)) dut(
		.clk(clk),
		.reset(reset),
		.MTimerInt(MTimerInt),
		.MExtInt(MExtInt),
		.SExtInt(SExtInt),
		.MSwInt(MSwInt),
		.MTIME_CLINT(MTIME_CLINT),
		.HRDATA(HRDATA),
		.HREADY(HREADY),
		.HRESP(HRESP),
		.HCLK(HCLK),
		.HRESETn(HRESETn),
		.HADDR(HADDR),
		.HWDATA(HWDATA),
		.HWSTRB(HWSTRB),
		.HWRITE(HWRITE),
		.HSIZE(HSIZE),
		.HBURST(HBURST),
		.HPROT(HPROT),
		.HTRANS(HTRANS),
		.HMASTLOCK(HMASTLOCK),
		.ExternalStall(ExternalStall)
	);
endmodule
module cache (
	clk,
	reset,
	Stall,
	FlushStage,
	CacheRW,
	FlushCache,
	InvalidateCache,
	CMOpM,
	NextSet,
	PAdr,
	ByteMask,
	WriteData,
	CacheCommitted,
	CacheStall,
	ReadDataWord,
	CacheMiss,
	CacheAccess,
	SelHPTW,
	CacheBusAck,
	SelBusBeat,
	BeatCount,
	FetchBuffer,
	CacheBusRW,
	CacheBusAdr
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter PA_BITS = 0;
	parameter LINELEN = 0;
	parameter NUMSETS = 0;
	parameter NUMWAYS = 4;
	parameter LOGBWPL = 0;
	parameter WORDLEN = 0;
	parameter MUXINTERVAL = 0;
	parameter READ_ONLY_CACHE = 0;
	input wire clk;
	input wire reset;
	input wire Stall;
	input wire FlushStage;
	input wire [1:0] CacheRW;
	input wire FlushCache;
	input wire InvalidateCache;
	input wire [3:0] CMOpM;
	input wire [11:0] NextSet;
	input wire [PA_BITS - 1:0] PAdr;
	input wire [(WORDLEN - 1) / 8:0] ByteMask;
	input wire [WORDLEN - 1:0] WriteData;
	output wire CacheCommitted;
	output wire CacheStall;
	output wire [WORDLEN - 1:0] ReadDataWord;
	output wire CacheMiss;
	output wire CacheAccess;
	input wire SelHPTW;
	input wire CacheBusAck;
	input wire SelBusBeat;
	input wire [LOGBWPL - 1:0] BeatCount;
	input wire [LINELEN - 1:0] FetchBuffer;
	output wire [1:0] CacheBusRW;
	output wire [PA_BITS - 1:0] CacheBusAdr;
	localparam LINEBYTELEN = LINELEN / 8;
	localparam OFFSETLEN = $clog2(LINEBYTELEN);
	localparam SETLEN = $clog2(NUMSETS);
	localparam SETTOP = SETLEN + OFFSETLEN;
	localparam TAGLEN = PA_BITS - SETTOP;
	localparam FLUSHADRTHRESHOLD = NUMSETS - 1;
	wire SelAdrData;
	wire SelAdrTag;
	wire [1:0] AdrSelMuxSelData;
	wire [1:0] AdrSelMuxSelTag;
	wire [1:0] AdrSelMuxSelLRU;
	wire [SETLEN - 1:0] CacheSetData;
	wire [SETLEN - 1:0] CacheSetTag;
	wire [SETLEN - 1:0] CacheSetLRU;
	wire [LINELEN - 1:0] LineWriteData;
	wire ClearDirty;
	wire SetDirty;
	wire SetValid;
	wire ClearValid;
	wire [(NUMWAYS * LINELEN) - 1:0] ReadDataLineWay;
	wire [NUMWAYS - 1:0] HitWay;
	wire [NUMWAYS - 1:0] ValidWay;
	wire Hit;
	wire [NUMWAYS - 1:0] VictimWay;
	wire [NUMWAYS - 1:0] DirtyWay;
	wire [NUMWAYS - 1:0] HitDirtyWay;
	wire LineDirty;
	wire HitLineDirty;
	wire [(NUMWAYS * TAGLEN) - 1:0] TagWay;
	wire [TAGLEN - 1:0] Tag;
	wire [SETLEN - 1:0] FlushAdr;
	wire FlushAdrCntEn;
	wire FlushCntRst;
	wire FlushAdrFlag;
	wire FlushWayFlag;
	wire [NUMWAYS - 1:0] FlushWay;
	wire [NUMWAYS - 1:0] NextFlushWay;
	wire FlushWayCntEn;
	wire SelWriteback;
	wire LRUWriteEn;
	wire [LINELEN - 1:0] ReadDataLine;
	wire [LINELEN - 1:0] ReadDataLineCache;
	wire SelFetchBuffer;
	wire CacheEn;
	wire SelVictim;
	wire [(LINELEN / 8) - 1:0] LineByteMask;
	wire [($clog2(LINELEN / 8) - $clog2(MUXINTERVAL / 8)) - 1:0] WordOffsetAddr;
	genvar _gv_index_1;
	assign AdrSelMuxSelData = {FlushCache, (SelAdrData | SelHPTW) & ~((READ_ONLY_CACHE == 1) & FlushStage)};
	mux3 #(.WIDTH(SETLEN)) AdrSelMuxData(
		.d0(NextSet[SETTOP - 1:OFFSETLEN]),
		.d1(PAdr[SETTOP - 1:OFFSETLEN]),
		.d2(FlushAdr),
		.s(AdrSelMuxSelData),
		.y(CacheSetData)
	);
	assign AdrSelMuxSelTag = {FlushCache, (SelAdrTag | SelHPTW) & ~((READ_ONLY_CACHE == 1) & FlushStage)};
	mux3 #(.WIDTH(SETLEN)) AdrSelMuxTag(
		.d0(NextSet[SETTOP - 1:OFFSETLEN]),
		.d1(PAdr[SETTOP - 1:OFFSETLEN]),
		.d2(FlushAdr),
		.s(AdrSelMuxSelTag),
		.y(CacheSetTag)
	);
	assign AdrSelMuxSelLRU = {FlushCache, ((SelAdrTag | SelHPTW) | Stall) & ~((READ_ONLY_CACHE == 1) & FlushStage)};
	mux3 #(.WIDTH(SETLEN)) AdrSelMuxLRU(
		.d0(NextSet[SETTOP - 1:OFFSETLEN]),
		.d1(PAdr[SETTOP - 1:OFFSETLEN]),
		.d2(FlushAdr),
		.s(AdrSelMuxSelLRU),
		.y(CacheSetLRU)
	);
	cacheway #(
		.P(P),
		.PA_BITS(PA_BITS),
		.NUMSETS(NUMSETS),
		.LINELEN(LINELEN),
		.TAGLEN(TAGLEN),
		.OFFSETLEN(OFFSETLEN),
		.INDEXLEN(SETLEN),
		.READ_ONLY_CACHE(READ_ONLY_CACHE)
	) CacheWays[NUMWAYS - 1:0](
		.clk(clk),
		.reset(reset),
		.CacheEn(CacheEn),
		.CacheSetData(CacheSetData),
		.CacheSetTag(CacheSetTag),
		.PAdr(PAdr),
		.LineWriteData(LineWriteData),
		.LineByteMask(LineByteMask),
		.SelVictim(SelVictim),
		.SetValid(SetValid),
		.ClearValid(ClearValid),
		.SetDirty(SetDirty),
		.ClearDirty(ClearDirty),
		.VictimWay(VictimWay),
		.FlushWay(FlushWay),
		.FlushCache(FlushCache),
		.ReadDataLineWay(ReadDataLineWay),
		.HitWay(HitWay),
		.ValidWay(ValidWay),
		.DirtyWay(DirtyWay),
		.HitDirtyWay(HitDirtyWay),
		.TagWay(TagWay),
		.FlushStage(FlushStage),
		.InvalidateCache(InvalidateCache)
	);
	generate
		if (NUMWAYS > 1) begin : vict
			cacheLRU #(
				.NUMWAYS(NUMWAYS),
				.SETLEN(SETLEN),
				.NUMSETS(NUMSETS)
			) cacheLRU(
				.clk(clk),
				.reset(reset),
				.FlushStage(FlushStage),
				.CacheEn(CacheEn),
				.HitWay(HitWay),
				.ValidWay(ValidWay),
				.VictimWay(VictimWay),
				.CacheSetLRU(CacheSetLRU),
				.LRUWriteEn(LRUWriteEn),
				.SetValid(SetValid),
				.PAdr(PAdr[SETTOP - 1:OFFSETLEN]),
				.InvalidateCache(InvalidateCache)
			);
		end
		else begin : genblk1
			assign VictimWay = 1'b1;
		end
	endgenerate
	assign Hit = |HitWay;
	assign LineDirty = |DirtyWay;
	assign HitLineDirty = |HitDirtyWay;
	or_rows #(
		.ROWS(NUMWAYS),
		.COLS(LINELEN)
	) ReadDataAOMux(
		.a(ReadDataLineWay),
		.y(ReadDataLineCache)
	);
	or_rows #(
		.ROWS(NUMWAYS),
		.COLS(TAGLEN)
	) TagAOMux(
		.a(TagWay),
		.y(Tag)
	);
	generate
		if (!READ_ONLY_CACHE) begin : genblk2
			mux2 #(.WIDTH(LOGBWPL)) WordAdrrMux(
				.d0(PAdr[$clog2(LINELEN / 8) - 1:$clog2(MUXINTERVAL / 8)]),
				.d1(BeatCount),
				.s(SelBusBeat),
				.y(WordOffsetAddr)
			);
		end
		else begin : genblk2
			assign WordOffsetAddr = PAdr[$clog2(LINELEN / 8) - 1:$clog2(MUXINTERVAL / 8)];
		end
	endgenerate
	mux2 #(.WIDTH(LINELEN)) EarlyReturnMux(
		.d0(ReadDataLineCache),
		.d1(FetchBuffer),
		.s(SelFetchBuffer),
		.y(ReadDataLine)
	);
	subcachelineread #(
		.LINELEN(LINELEN),
		.WORDLEN(WORDLEN),
		.MUXINTERVAL(MUXINTERVAL)
	) subcachelineread(
		.PAdr(WordOffsetAddr),
		.ReadDataLine(ReadDataLine),
		.ReadDataWord(ReadDataWord)
	);
	mux3 #(.WIDTH(PA_BITS)) CacheBusAdrMux(
		.d0({PAdr[PA_BITS - 1:OFFSETLEN], {OFFSETLEN {1'b0}}}),
		.d1({Tag, PAdr[SETTOP - 1:OFFSETLEN], {OFFSETLEN {1'b0}}}),
		.d2({Tag, FlushAdr, {OFFSETLEN {1'b0}}}),
		.s({FlushCache, SelWriteback}),
		.y(CacheBusAdr)
	);
	generate
		if (!READ_ONLY_CACHE) begin : WriteSelLogic
			wire [(LINELEN / 8) - 1:0] DemuxedByteMask;
			wire [(LINELEN / 8) - 1:0] FetchBufferByteSel;
			wire [(LINELEN / 8) - 1:0] BlankByteMask;
			assign BlankByteMask[(WORDLEN / 8) - 1:0] = ByteMask;
			assign BlankByteMask[(LINELEN / 8) - 1:WORDLEN / 8] = 0;
			assign DemuxedByteMask = BlankByteMask << ((MUXINTERVAL / 8) * WordOffsetAddr);
			assign FetchBufferByteSel = (SetDirty ? ~DemuxedByteMask : {LINELEN / 8 {1'sb1}});
			for (_gv_index_1 = 0; _gv_index_1 < (LINELEN / 8); _gv_index_1 = _gv_index_1 + 1) begin : genblk1
				localparam index = _gv_index_1;
				mux2 #(.WIDTH(8)) WriteDataMux(
					.d0(WriteData[((8 * index) % WORDLEN) + 7:(8 * index) % WORDLEN]),
					.d1(FetchBuffer[(8 * index) + 7:8 * index]),
					.s(FetchBufferByteSel[index] & ~CMOpM[3]),
					.y(LineWriteData[(8 * index) + 7:8 * index])
				);
			end
			assign LineByteMask = (SetDirty ? DemuxedByteMask : {LINELEN / 8 {1'sb1}});
		end
		else begin : WriteSelLogic
			assign LineWriteData = FetchBuffer;
			assign LineByteMask = 1'sb1;
		end
		if (!READ_ONLY_CACHE) begin : flushlogic
			wire ResetOrFlushCntRst;
			wire [SETLEN - 1:0] NextFlushAdr;
			wire [SETLEN - 1:0] FlushAdrP1;
			assign ResetOrFlushCntRst = reset | FlushCntRst;
			flopenr #(.WIDTH(SETLEN)) FlushAdrReg(
				.clk(clk),
				.reset(ResetOrFlushCntRst),
				.en(FlushAdrCntEn),
				.d(FlushAdrP1),
				.q(NextFlushAdr)
			);
			mux2 #(.WIDTH(SETLEN)) FlushAdrMux(
				.d0(NextFlushAdr),
				.d1(FlushAdrP1),
				.s(FlushAdrCntEn),
				.y(FlushAdr)
			);
			assign FlushAdrP1 = NextFlushAdr + 1'b1;
			assign FlushAdrFlag = NextFlushAdr == FLUSHADRTHRESHOLD[SETLEN - 1:0];
			flopenl #(.WIDTH(NUMWAYS)) FlushWayReg(
				.clk(clk),
				.load(FlushWayCntEn),
				.en(ResetOrFlushCntRst),
				.d({{NUMWAYS - 1 {1'b0}}, 1'b1}),
				.val(NextFlushWay),
				.q(FlushWay)
			);
			if (NUMWAYS > 1) begin : genblk1
				assign NextFlushWay = {FlushWay[NUMWAYS - 2:0], FlushWay[NUMWAYS - 1]};
			end
			else begin : genblk1
				assign NextFlushWay = FlushWay[NUMWAYS - 1];
			end
			assign FlushWayFlag = FlushWay[NUMWAYS - 1];
		end
		else begin : flushlogic
			assign FlushWay = 1'sb0;
			assign FlushWayFlag = 1'b0;
			assign FlushAdrFlag = 1'b0;
			assign FlushAdr = 1'sb0;
		end
	endgenerate
	cachefsm #(.READ_ONLY_CACHE(READ_ONLY_CACHE)) cachefsm(
		.clk(clk),
		.reset(reset),
		.CacheBusRW(CacheBusRW),
		.CacheBusAck(CacheBusAck),
		.FlushStage(FlushStage),
		.CacheRW(CacheRW),
		.Stall(Stall),
		.Hit(Hit),
		.LineDirty(LineDirty),
		.HitLineDirty(HitLineDirty),
		.CacheStall(CacheStall),
		.CacheCommitted(CacheCommitted),
		.CacheMiss(CacheMiss),
		.CacheAccess(CacheAccess),
		.SelAdrData(SelAdrData),
		.SelAdrTag(SelAdrTag),
		.SelVictim(SelVictim),
		.ClearDirty(ClearDirty),
		.SetDirty(SetDirty),
		.SetValid(SetValid),
		.ClearValid(ClearValid),
		.SelWriteback(SelWriteback),
		.FlushAdrCntEn(FlushAdrCntEn),
		.FlushWayCntEn(FlushWayCntEn),
		.FlushCntRst(FlushCntRst),
		.FlushAdrFlag(FlushAdrFlag),
		.FlushWayFlag(FlushWayFlag),
		.FlushCache(FlushCache),
		.SelFetchBuffer(SelFetchBuffer),
		.InvalidateCache(InvalidateCache),
		.CMOpM(CMOpM),
		.CacheEn(CacheEn),
		.LRUWriteEn(LRUWriteEn)
	);
endmodule
module cachefsm (
	clk,
	reset,
	Stall,
	FlushStage,
	CacheCommitted,
	CacheStall,
	CacheRW,
	FlushCache,
	InvalidateCache,
	CMOpM,
	CacheBusAck,
	CacheBusRW,
	CacheMiss,
	CacheAccess,
	Hit,
	LineDirty,
	HitLineDirty,
	FlushAdrFlag,
	FlushWayFlag,
	SelAdrData,
	SelAdrTag,
	SetValid,
	ClearValid,
	SetDirty,
	ClearDirty,
	SelWriteback,
	LRUWriteEn,
	SelVictim,
	FlushAdrCntEn,
	FlushWayCntEn,
	FlushCntRst,
	SelFetchBuffer,
	CacheEn
);
	reg _sv2v_0;
	parameter READ_ONLY_CACHE = 0;
	input wire clk;
	input wire reset;
	input wire Stall;
	input wire FlushStage;
	output wire CacheCommitted;
	output wire CacheStall;
	input wire [1:0] CacheRW;
	input wire FlushCache;
	input wire InvalidateCache;
	input wire [3:0] CMOpM;
	input wire CacheBusAck;
	output wire [1:0] CacheBusRW;
	output wire CacheMiss;
	output wire CacheAccess;
	input wire Hit;
	input wire LineDirty;
	input wire HitLineDirty;
	input wire FlushAdrFlag;
	input wire FlushWayFlag;
	output wire SelAdrData;
	output wire SelAdrTag;
	output wire SetValid;
	output wire ClearValid;
	output wire SetDirty;
	output wire ClearDirty;
	output wire SelWriteback;
	output wire LRUWriteEn;
	output wire SelVictim;
	output wire FlushAdrCntEn;
	output wire FlushWayCntEn;
	output wire FlushCntRst;
	output wire SelFetchBuffer;
	output wire CacheEn;
	wire resetDelay;
	wire AnyUpdateHit;
	wire AnyHit;
	wire AnyMiss;
	wire FlushFlag;
	wire CMOWriteback;
	wire CMOZeroNoEviction;
	wire StallConditions;
	reg [3:0] CurrState;
	reg [3:0] NextState;
	assign AnyMiss = ((CacheRW[0] | CacheRW[1]) & ~Hit) & ~InvalidateCache;
	assign AnyUpdateHit = CacheRW[0] & Hit;
	assign AnyHit = AnyUpdateHit | (CacheRW[1] & Hit);
	assign CMOZeroNoEviction = CMOpM[3] & ~LineDirty;
	assign CMOWriteback = (((CMOpM[1] | CMOpM[2]) & Hit) & HitLineDirty) | (CMOpM[3] & LineDirty);
	assign FlushFlag = FlushAdrFlag & FlushWayFlag;
	assign CacheAccess = |CacheRW & ((((CurrState == 4'd0) & ~Stall) & ~FlushStage) | (((CurrState == 4'd4) & ~Stall) & ~FlushStage));
	assign CacheMiss = ((CurrState == 4'd4) & ~Stall) & ~FlushStage;
	flop #(.WIDTH(1)) resetDelayReg(
		.clk(clk),
		.d(reset),
		.q(resetDelay)
	);
	always @(posedge clk)
		if (reset | FlushStage)
			CurrState <= 4'd0;
		else
			CurrState <= NextState;
	always @(*) begin
		if (_sv2v_0)
			;
		NextState = 4'd0;
		case (CurrState)
			4'd0:
				if (InvalidateCache)
					NextState = 4'd0;
				else if (FlushCache & ~READ_ONLY_CACHE)
					NextState = 4'd5;
				else if (AnyMiss & (READ_ONLY_CACHE | ~LineDirty))
					NextState = 4'd1;
				else if ((AnyMiss | CMOWriteback) & ~READ_ONLY_CACHE)
					NextState = 4'd2;
				else
					NextState = 4'd0;
			4'd1:
				if (CacheBusAck)
					NextState = 4'd3;
				else
					NextState = 4'd1;
			4'd3: NextState = 4'd4;
			4'd4:
				if (Stall)
					NextState = 4'd4;
				else
					NextState = 4'd0;
			4'd2:
				if (CacheBusAck & ~(|CMOpM[3:1]))
					NextState = 4'd1;
				else if (CacheBusAck)
					NextState = 4'd4;
				else
					NextState = 4'd2;
			4'd5:
				if (LineDirty)
					NextState = 4'd6;
				else if (FlushFlag)
					NextState = 4'd4;
				else
					NextState = 4'd5;
			4'd6:
				if (CacheBusAck & ~FlushFlag)
					NextState = 4'd5;
				else if (CacheBusAck)
					NextState = 4'd4;
				else
					NextState = 4'd6;
			default: NextState = 4'd0;
		endcase
	end
	assign CacheCommitted = (CurrState != 4'd0) & ~(READ_ONLY_CACHE & (CurrState == 4'd4));
	assign StallConditions = (FlushCache | AnyMiss) | CMOWriteback;
	assign CacheStall = ((((((CurrState == 4'd0) & StallConditions) | (CurrState == 4'd1)) | (CurrState == 4'd2)) | (CurrState == 4'd3)) | (CurrState == 4'd5)) | (CurrState == 4'd6);
	assign SetValid = ((CurrState == 4'd3) | ((CurrState == 4'd0) & CMOZeroNoEviction)) | (((CurrState == 4'd2) & CacheBusAck) & CMOpM[3]);
	assign ClearValid = ((CurrState == 4'd0) & (CMOpM[0] | (CMOpM[2] & ~HitLineDirty))) | (((CurrState == 4'd2) & CMOpM[2]) & CacheBusAck);
	assign LRUWriteEn = ((((CurrState == 4'd0) & (AnyHit | CMOZeroNoEviction)) | (CurrState == 4'd3)) & ~FlushStage) | (((CurrState == 4'd2) & CMOpM[3]) & CacheBusAck);
	assign SetDirty = (((CurrState == 4'd0) & (AnyUpdateHit | CMOZeroNoEviction)) | ((CurrState == 4'd3) & CacheRW[0])) | ((CurrState == 4'd2) & (CMOpM[3] & CacheBusAck));
	assign ClearDirty = (((CurrState == 4'd3) & ~CacheRW[0]) | ((CurrState == 4'd5) & LineDirty)) | (((CurrState == 4'd2) & (CMOpM[1] | CMOpM[2])) & CacheBusAck);
	assign SelVictim = (((CurrState == 4'd2) & ((~CacheBusAck & ~(CMOpM[1] | CMOpM[2])) | (CacheBusAck & CMOpM[3]))) | ((CurrState == 4'd0) & ((AnyMiss & LineDirty) | (CMOZeroNoEviction & ~Hit)))) | (CurrState == 4'd3);
	assign SelWriteback = ((CurrState == 4'd2) & ((CMOpM[1] | CMOpM[2]) | ~CacheBusAck)) | (((CurrState == 4'd0) & AnyMiss) & LineDirty);
	assign FlushAdrCntEn = (((CurrState == 4'd6) & FlushWayFlag) & CacheBusAck) | (((CurrState == 4'd5) & FlushWayFlag) & ~LineDirty);
	assign FlushWayCntEn = ((CurrState == 4'd5) & ~LineDirty) | ((CurrState == 4'd6) & CacheBusAck);
	assign FlushCntRst = (((CurrState == 4'd5) & FlushFlag) & ~LineDirty) | (((CurrState == 4'd6) & FlushFlag) & CacheBusAck);
	assign CacheBusRW[1] = ((((CurrState == 4'd0) & AnyMiss) & ~LineDirty) | ((CurrState == 4'd1) & ~CacheBusAck)) | (((CurrState == 4'd2) & CacheBusAck) & ~(|CMOpM));
	wire LoadMiss;
	assign LoadMiss = (CacheRW[1] & ~Hit) & ~InvalidateCache;
	assign CacheBusRW[0] = (((((CurrState == 4'd0) & LoadMiss) & LineDirty) | ((CurrState == 4'd2) & ~CacheBusAck)) | ((CurrState == 4'd6) & ~CacheBusAck)) | (((CurrState == 4'd2) & (CMOpM[1] | CMOpM[2])) & ~CacheBusAck);
	assign SelAdrData = (((((CurrState == 4'd0) & ((CacheRW[0] | AnyMiss) | (|CMOpM))) | (CurrState == 4'd1)) | (CurrState == 4'd2)) | (CurrState == 4'd3)) | resetDelay;
	assign SelAdrTag = (((((CurrState == 4'd0) & (AnyMiss | (|CMOpM))) | (CurrState == 4'd1)) | (CurrState == 4'd2)) | (CurrState == 4'd3)) | resetDelay;
	assign SelFetchBuffer = (CurrState == 4'd3) | (CurrState == 4'd4);
	assign CacheEn = (((~Stall | StallConditions) | (CurrState != 4'd0)) | reset) | InvalidateCache;
	initial _sv2v_0 = 0;
endmodule
module cacheway (
	clk,
	reset,
	FlushStage,
	CacheEn,
	CacheSetData,
	CacheSetTag,
	PAdr,
	LineWriteData,
	SetValid,
	ClearValid,
	SetDirty,
	SelVictim,
	ClearDirty,
	FlushCache,
	VictimWay,
	FlushWay,
	InvalidateCache,
	LineByteMask,
	ReadDataLineWay,
	HitWay,
	ValidWay,
	HitDirtyWay,
	DirtyWay,
	TagWay
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter PA_BITS = 0;
	parameter NUMSETS = 512;
	parameter LINELEN = 256;
	parameter TAGLEN = 26;
	parameter OFFSETLEN = 5;
	parameter INDEXLEN = 9;
	parameter READ_ONLY_CACHE = 0;
	input wire clk;
	input wire reset;
	input wire FlushStage;
	input wire CacheEn;
	input wire [$clog2(NUMSETS) - 1:0] CacheSetData;
	input wire [$clog2(NUMSETS) - 1:0] CacheSetTag;
	input wire [PA_BITS - 1:0] PAdr;
	input wire [LINELEN - 1:0] LineWriteData;
	input wire SetValid;
	input wire ClearValid;
	input wire SetDirty;
	input wire SelVictim;
	input wire ClearDirty;
	input wire FlushCache;
	input wire VictimWay;
	input wire FlushWay;
	input wire InvalidateCache;
	input wire [(LINELEN / 8) - 1:0] LineByteMask;
	output wire [LINELEN - 1:0] ReadDataLineWay;
	output wire HitWay;
	output reg ValidWay;
	output wire HitDirtyWay;
	output wire DirtyWay;
	output wire [TAGLEN - 1:0] TagWay;
	reg [NUMSETS - 1:0] ValidBits;
	reg [NUMSETS - 1:0] DirtyBits;
	wire [LINELEN - 1:0] ReadDataLine;
	wire [TAGLEN - 1:0] ReadTag;
	reg Dirty;
	wire SelecteDirty;
	wire SelectedWriteWordEn;
	wire [(LINELEN / 8) - 1:0] FinalByteMask;
	wire SetValidEN;
	wire ClearValidEN;
	wire SetValidWay;
	wire ClearValidWay;
	wire SetDirtyWay;
	wire ClearDirtyWay;
	wire SelectedWay;
	wire InvalidateCacheDelay;
	generate
		if (!READ_ONLY_CACHE) begin : flushlogic
			mux2 #(.WIDTH(1)) seltagmux(
				.d0(VictimWay),
				.d1(FlushWay),
				.s(FlushCache),
				.y(SelecteDirty)
			);
			mux3 #(.WIDTH(1)) selectedmux(
				.d0(HitWay),
				.d1(FlushWay),
				.d2(VictimWay),
				.s({SelVictim, FlushCache}),
				.y(SelectedWay)
			);
		end
		else begin : flushlogic
			assign SelecteDirty = VictimWay;
			mux2 #(.WIDTH(1)) selectedwaymux(
				.d0(HitWay),
				.d1(SelecteDirty),
				.s(SelVictim),
				.y(SelectedWay)
			);
		end
	endgenerate
	assign SetValidWay = SetValid & SelectedWay;
	assign ClearValidWay = ClearValid & SelectedWay;
	assign SetDirtyWay = SetDirty & SelectedWay;
	assign ClearDirtyWay = ClearDirty & SelectedWay;
	assign SelectedWriteWordEn = (SetValidWay | SetDirtyWay) & ~FlushStage;
	assign SetValidEN = SetValidWay & ~FlushStage;
	assign ClearValidEN = ClearValidWay & ~FlushStage;
	assign FinalByteMask = (SetValidWay ? {LINELEN / 8 {1'sb1}} : LineByteMask);
	ram1p1rwe #(
		.USE_SRAM(P[1743]),
		.DEPTH(NUMSETS),
		.WIDTH(TAGLEN)
	) CacheTagMem(
		.clk(clk),
		.ce(CacheEn),
		.addr(CacheSetTag),
		.dout(ReadTag),
		.din(PAdr[PA_BITS - 1:OFFSETLEN + INDEXLEN]),
		.we(SetValidEN)
	);
	assign TagWay = (SelectedWay ? ReadTag : 0);
	assign HitDirtyWay = Dirty & ValidWay;
	assign DirtyWay = SelecteDirty & HitDirtyWay;
	assign HitWay = (ValidWay & (ReadTag == PAdr[PA_BITS - 1:OFFSETLEN + INDEXLEN])) & ~InvalidateCacheDelay;
	flop #(.WIDTH(1)) InvalidateCacheReg(
		.clk(clk),
		.d(InvalidateCache),
		.q(InvalidateCacheDelay)
	);
	genvar _gv_words_1;
	localparam NUMSRAM = LINELEN / $signed(P[3793-:32]);
	localparam SRAMLENINBYTES = $signed(P[3793-:32]) / 8;
	generate
		for (_gv_words_1 = 0; _gv_words_1 < NUMSRAM; _gv_words_1 = _gv_words_1 + 1) begin : word
			localparam words = _gv_words_1;
			if (READ_ONLY_CACHE) begin : wordram
				ram1p1rwe #(
					.USE_SRAM(P[1743]),
					.DEPTH(NUMSETS),
					.WIDTH($signed(P[3793-:32]))
				) CacheDataMem(
					.clk(clk),
					.ce(CacheEn),
					.addr(CacheSetData),
					.dout(ReadDataLine[($signed(P[3793-:32]) * (words + 1)) - 1:$signed(P[3793-:32]) * words]),
					.din(LineWriteData[($signed(P[3793-:32]) * (words + 1)) - 1:$signed(P[3793-:32]) * words]),
					.we(SelectedWriteWordEn)
				);
			end
			else begin : wordram
				ram1p1rwbe #(
					.USE_SRAM(P[1743]),
					.DEPTH(NUMSETS),
					.WIDTH($signed(P[3793-:32]))
				) CacheDataMem(
					.clk(clk),
					.ce(CacheEn),
					.addr(CacheSetData),
					.dout(ReadDataLine[($signed(P[3793-:32]) * (words + 1)) - 1:$signed(P[3793-:32]) * words]),
					.din(LineWriteData[($signed(P[3793-:32]) * (words + 1)) - 1:$signed(P[3793-:32]) * words]),
					.we(SelectedWriteWordEn),
					.bwe(FinalByteMask[(SRAMLENINBYTES * (words + 1)) - 1:SRAMLENINBYTES * words])
				);
			end
		end
	endgenerate
	assign ReadDataLineWay = (SelectedWay ? ReadDataLine : {LINELEN {1'sb0}});
	always @(posedge clk) begin
		if (reset)
			ValidBits <= 1'sb0;
		if (CacheEn) begin
			ValidWay <= ValidBits[CacheSetTag];
			if (InvalidateCache)
				ValidBits <= 1'sb0;
			else if (SetValidEN)
				ValidBits[CacheSetData] <= SetValidWay;
			else if (ClearValidEN)
				ValidBits[CacheSetData] <= 1'sb0;
		end
	end
	generate
		if (!READ_ONLY_CACHE) begin : dirty
			always @(posedge clk)
				if (CacheEn) begin
					Dirty <= DirtyBits[CacheSetTag];
					if ((SetDirtyWay | ClearDirtyWay) & ~FlushStage) begin
						DirtyBits[CacheSetData] <= SetDirtyWay;
						if (CacheSetData == CacheSetTag)
							Dirty <= SetDirtyWay;
						else
							Dirty <= DirtyBits[CacheSetTag];
					end
				end
		end
		else begin : genblk3
			wire [1:1] sv2v_tmp_ABFB2;
			assign sv2v_tmp_ABFB2 = 1'b0;
			always @(*) Dirty = sv2v_tmp_ABFB2;
		end
	endgenerate
endmodule
module subcachelineread (
	PAdr,
	ReadDataLine,
	ReadDataWord
);
	parameter LINELEN = 0;
	parameter WORDLEN = 0;
	parameter MUXINTERVAL = 0;
	input wire [($clog2(LINELEN / 8) - $clog2(MUXINTERVAL / 8)) - 1:0] PAdr;
	input wire [LINELEN - 1:0] ReadDataLine;
	output wire [WORDLEN - 1:0] ReadDataWord;
	localparam WORDSPERLINE = LINELEN / MUXINTERVAL;
	localparam PADLEN = WORDLEN - MUXINTERVAL;
	wire [(LINELEN + (WORDLEN - MUXINTERVAL)) - 1:0] ReadDataLinePad;
	wire [WORDLEN - 1:0] ReadDataLineSets [(LINELEN / MUXINTERVAL) - 1:0];
	generate
		if (PADLEN > 0) begin : genblk1
			assign ReadDataLinePad = {{PADLEN {1'b0}}, ReadDataLine};
		end
		else begin : genblk1
			assign ReadDataLinePad = ReadDataLine;
		end
	endgenerate
	genvar _gv_index_2;
	generate
		for (_gv_index_2 = 0; _gv_index_2 < WORDSPERLINE; _gv_index_2 = _gv_index_2 + 1) begin : readdatalinesetsmux
			localparam index = _gv_index_2;
			assign ReadDataLineSets[index] = ReadDataLinePad[((index * MUXINTERVAL) + WORDLEN) - 1:index * MUXINTERVAL];
		end
	endgenerate
	assign ReadDataWord = ReadDataLineSets[PAdr];
endmodule
module cacheLRU (
	clk,
	reset,
	FlushStage,
	CacheEn,
	HitWay,
	ValidWay,
	CacheSetLRU,
	PAdr,
	LRUWriteEn,
	SetValid,
	InvalidateCache,
	VictimWay
);
	parameter NUMWAYS = 4;
	parameter SETLEN = 9;
	parameter NUMSETS = 128;
	input wire clk;
	input wire reset;
	input wire FlushStage;
	input wire CacheEn;
	input wire [NUMWAYS - 1:0] HitWay;
	input wire [NUMWAYS - 1:0] ValidWay;
	input wire [SETLEN - 1:0] CacheSetLRU;
	input wire [SETLEN - 1:0] PAdr;
	input wire LRUWriteEn;
	input wire SetValid;
	input wire InvalidateCache;
	output wire [NUMWAYS - 1:0] VictimWay;
	localparam LOGNUMWAYS = $clog2(NUMWAYS);
	reg [NUMWAYS - 2:0] LRUMemory [NUMSETS - 1:0];
	wire [NUMWAYS - 2:0] CurrLRU;
	wire [NUMWAYS - 2:0] NextLRU;
	wire [NUMWAYS - 2:0] ReadLRU;
	wire [NUMWAYS - 2:0] BypassedLRU;
	wire [LOGNUMWAYS - 1:0] HitWayEncoded;
	wire [LOGNUMWAYS - 1:0] Way;
	wire [NUMWAYS - 2:0] WayExpanded;
	wire AllValid;
	wire ForwardLRU;
	genvar _gv_row_1;
	wire [NUMWAYS - 2:0] LRUUpdate;
	wire [LOGNUMWAYS - 1:0] Intermediate [NUMWAYS - 2:0];
	wire [NUMWAYS - 1:0] FirstZero;
	wire [LOGNUMWAYS - 1:0] FirstZeroWay;
	wire [LOGNUMWAYS - 1:0] VictimWayEnc;
	binencoder #(.N(NUMWAYS)) hitwayencoder(
		.A(HitWay),
		.Y(HitWayEncoded)
	);
	assign AllValid = &ValidWay;
	function integer log2;
		input integer value;
		reg signed [31:0] val;
		begin
			val = value;
			for (log2 = 0; val > 0; log2 = log2 + 1)
				val = val >> 1;
			log2 = log2;
		end
	endfunction
	mux2 #(.WIDTH(LOGNUMWAYS)) WayMuxEnc(
		.d0(HitWayEncoded),
		.d1(VictimWayEnc),
		.s(SetValid),
		.y(Way)
	);
	generate
		for (_gv_row_1 = 0; _gv_row_1 < LOGNUMWAYS; _gv_row_1 = _gv_row_1 + 1) begin : genblk1
			localparam row = _gv_row_1;
			localparam integer DuplicationFactor = 2 ** ((LOGNUMWAYS - row) - 1);
			localparam StartIndex = ((NUMWAYS - 2) - DuplicationFactor) + 1;
			localparam EndIndex = ((NUMWAYS - 2) - (2 * DuplicationFactor)) + 2;
			assign WayExpanded[StartIndex:EndIndex] = {{DuplicationFactor} {Way[row]}};
		end
	endgenerate
	genvar _gv_node_1;
	assign LRUUpdate[NUMWAYS - 2] = 1'sb1;
	generate
		for (_gv_node_1 = NUMWAYS - 2; _gv_node_1 >= (NUMWAYS / 2); _gv_node_1 = _gv_node_1 - 1) begin : enables
			localparam node = _gv_node_1;
			localparam ctr = (NUMWAYS - node) - 1;
			localparam ctr_depth = log2(ctr);
			localparam lchild = node - ctr;
			localparam rchild = lchild - 1;
			localparam r = LOGNUMWAYS - ctr_depth;
			if (node == (NUMWAYS - 2)) begin : genblk1
				assign LRUUpdate[lchild] = ~Way[r];
				assign LRUUpdate[rchild] = Way[r];
			end
			else begin : genblk1
				assign LRUUpdate[lchild] = LRUUpdate[node] & ~Way[r];
				assign LRUUpdate[rchild] = LRUUpdate[node] & Way[r];
			end
		end
	endgenerate
	assign NextLRU[NUMWAYS - 2] = ~WayExpanded[NUMWAYS - 2];
	generate
		if (NUMWAYS > 2) begin : genblk3
			mux2 #(.WIDTH(1)) LRUMuxes[NUMWAYS - 3:0](
				.d0(CurrLRU[NUMWAYS - 3:0]),
				.d1(~WayExpanded[NUMWAYS - 3:0]),
				.s(LRUUpdate[NUMWAYS - 3:0]),
				.y(NextLRU[NUMWAYS - 3:0])
			);
		end
		for (_gv_node_1 = NUMWAYS - 2; _gv_node_1 >= (NUMWAYS / 2); _gv_node_1 = _gv_node_1 - 1) begin : genblk4
			localparam node = _gv_node_1;
			localparam t0 = (2 * node) - NUMWAYS;
			localparam t1 = t0 + 1;
			assign Intermediate[node] = (CurrLRU[node] ? Intermediate[t0] : Intermediate[t1]);
		end
		for (_gv_node_1 = (NUMWAYS >> 1) - 1; _gv_node_1 >= 0; _gv_node_1 = _gv_node_1 - 1) begin : genblk5
			localparam node = _gv_node_1;
			localparam int0 = (((NUMWAYS / 2) - 1) - node) * 2;
			localparam int1 = int0 + 1;
			assign Intermediate[node] = (CurrLRU[node] ? int1[LOGNUMWAYS - 1:0] : int0[LOGNUMWAYS - 1:0]);
		end
	endgenerate
	priorityonehot #(.N(NUMWAYS)) FirstZeroEncoder(
		.a(~ValidWay),
		.y(FirstZero)
	);
	binencoder #(.N(NUMWAYS)) FirstZeroWayEncoder(
		.A(FirstZero),
		.Y(FirstZeroWay)
	);
	mux2 #(.WIDTH(LOGNUMWAYS)) VictimMux(
		.d0(FirstZeroWay),
		.d1(Intermediate[NUMWAYS - 2]),
		.s(AllValid),
		.y(VictimWayEnc)
	);
	decoder #(.BINARY_BITS(LOGNUMWAYS)) decoder(
		.binary(VictimWayEnc),
		.onehot(VictimWay)
	);
	always @(posedge clk)
		if (reset | (InvalidateCache & ~FlushStage)) begin : sv2v_autoblock_1
			reg signed [31:0] set;
			for (set = 0; set < NUMSETS; set = set + 1)
				LRUMemory[set] <= 1'sb0;
		end
		else if (CacheEn & LRUWriteEn)
			LRUMemory[PAdr] <= NextLRU;
	assign ReadLRU = LRUMemory[CacheSetLRU];
	assign ForwardLRU = LRUWriteEn & (PAdr == CacheSetLRU);
	mux2 #(.WIDTH(NUMWAYS - 1)) ReadLRUmux(
		.d0(ReadLRU),
		.d1(NextLRU),
		.s(ForwardLRU),
		.y(BypassedLRU)
	);
	flop #(.WIDTH(NUMWAYS - 1)) CurrLRUReg(
		.clk(clk),
		.d(BypassedLRU),
		.q(CurrLRU)
	);
endmodule
module ahbcacheinterface (
	HCLK,
	HRESETn,
	HREADY,
	HTRANS,
	HWRITE,
	HSIZE,
	HBURST,
	HRDATA,
	HADDR,
	HWDATA,
	HWSTRB,
	CacheBusAdr,
	CacheReadDataWordM,
	CacheableOrFlushCacheM,
	Cacheable,
	CacheBusRW,
	CacheBusAck,
	FetchBuffer,
	BeatCount,
	SelBusBeat,
	PAdr,
	WriteDataM,
	BusRW,
	BusAtomic,
	Funct3,
	BusCMOZero,
	Stall,
	Flush,
	BusStall,
	BusCommitted
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter BEATSPERLINE = 0;
	parameter AHBWLOGBWPL = 0;
	parameter LINELEN = 0;
	parameter LLENPOVERAHBW = 0;
	parameter READ_ONLY_CACHE = 0;
	input wire HCLK;
	input wire HRESETn;
	input wire HREADY;
	output wire [1:0] HTRANS;
	output wire HWRITE;
	output wire [2:0] HSIZE;
	output wire [2:0] HBURST;
	input wire [$signed(P[4151-:32]) - 1:0] HRDATA;
	output wire [$signed(P[1640-:32]) - 1:0] HADDR;
	output wire [$signed(P[4151-:32]) - 1:0] HWDATA;
	output wire [($signed(P[4151-:32]) / 8) - 1:0] HWSTRB;
	input wire [$signed(P[1640-:32]) - 1:0] CacheBusAdr;
	input wire [$signed(P[383-:32]) - 1:0] CacheReadDataWordM;
	input wire CacheableOrFlushCacheM;
	input wire Cacheable;
	input wire [1:0] CacheBusRW;
	output wire CacheBusAck;
	output wire [LINELEN - 1:0] FetchBuffer;
	output wire [AHBWLOGBWPL - 1:0] BeatCount;
	output wire SelBusBeat;
	input wire [$signed(P[1640-:32]) - 1:0] PAdr;
	input wire [$signed(P[383-:32]) - 1:0] WriteDataM;
	input wire [1:0] BusRW;
	input wire BusAtomic;
	input wire [2:0] Funct3;
	input wire BusCMOZero;
	input wire Stall;
	input wire Flush;
	output wire BusStall;
	output wire BusCommitted;
	localparam BeatCountThreshold = BEATSPERLINE - 1;
	wire [$signed(P[1640-:32]) - 1:0] LocalHADDR;
	wire [AHBWLOGBWPL - 1:0] BeatCountDelayed;
	wire CaptureEn;
	wire [$signed(P[4151-:32]) - 1:0] PreHWDATA;
	wire [$signed(P[1640-:32]) - 1:0] PAdrZero;
	genvar _gv_index_3;
	generate
		for (_gv_index_3 = 0; _gv_index_3 < BEATSPERLINE; _gv_index_3 = _gv_index_3 + 1) begin : fetchbuffer
			localparam index = _gv_index_3;
			wire [BEATSPERLINE - 1:0] CaptureBeat;
			assign CaptureBeat[index] = CaptureEn & (index == BeatCountDelayed);
			flopen #(.WIDTH($signed(P[4151-:32]))) fb(
				.clk(HCLK),
				.en(CaptureBeat[index]),
				.d(HRDATA),
				.q(FetchBuffer[((index + 1) * $signed(P[4151-:32])) - 1:index * $signed(P[4151-:32])])
			);
		end
	endgenerate
	assign PAdrZero = (BusCMOZero ? {PAdr[$signed(P[1640-:32]) - 1:$clog2(LINELEN / 8)], {$clog2(LINELEN / 8) {1'b0}}} : PAdr);
	mux2 #(.WIDTH($signed(P[1640-:32]))) localadrmux(
		.d0(PAdrZero),
		.d1(CacheBusAdr),
		.s(Cacheable),
		.y(LocalHADDR)
	);
	assign HADDR = ({{$signed(P[1640-:32]) - AHBWLOGBWPL {1'b0}}, BeatCount} << $clog2($signed(P[4151-:32]) / 8)) + LocalHADDR;
	mux2 #(.WIDTH(3)) sizemux(
		.d0(Funct3),
		.d1(($signed(P[4151-:32]) == 32 ? 3'b010 : 3'b011)),
		.s(Cacheable | BusCMOZero),
		.y(HSIZE)
	);
	wire [$signed(P[4151-:32]) - 1:0] CacheReadDataWordAHB;
	generate
		if (LLENPOVERAHBW > 1) begin : genblk2
			wire [$signed(P[4151-:32]) - 1:0] AHBWordSets [LLENPOVERAHBW - 1:0];
			genvar _gv_index_4;
			for (_gv_index_4 = 0; _gv_index_4 < LLENPOVERAHBW; _gv_index_4 = _gv_index_4 + 1) begin : readdatalinesetsmux
				localparam index = _gv_index_4;
				assign AHBWordSets[index] = CacheReadDataWordM[((index * $signed(P[4151-:32])) + $signed(P[4151-:32])) - 1:index * $signed(P[4151-:32])];
			end
			assign CacheReadDataWordAHB = AHBWordSets[BeatCount[$clog2(LLENPOVERAHBW) - 1:0]];
		end
		else begin : genblk2
			assign CacheReadDataWordAHB = CacheReadDataWordM[$signed(P[4151-:32]) - 1:0];
		end
	endgenerate
	mux2 #(.WIDTH($signed(P[4151-:32]))) HWDATAMux(
		.d0(CacheReadDataWordAHB),
		.d1(WriteDataM[$signed(P[4151-:32]) - 1:0]),
		.s(~CacheableOrFlushCacheM),
		.y(PreHWDATA)
	);
	flopen #(.WIDTH($signed(P[4151-:32]))) wdreg(
		.clk(HCLK),
		.en(HREADY),
		.d(PreHWDATA),
		.q(HWDATA)
	);
	generate
		if (READ_ONLY_CACHE) begin : genblk3
			assign HWSTRB = 1'sb0;
		end
		else begin : genblk3
			wire [($signed(P[4151-:32]) / 8) - 1:0] BusByteMaskM;
			swbytemask #(.WORDLEN($signed(P[4151-:32]))) busswbytemask(
				.Size(HSIZE),
				.Adr(HADDR[$clog2($signed(P[4151-:32]) / 8) - 1:0]),
				.ByteMask(BusByteMaskM),
				.ByteMaskExtended()
			);
			flopen #(.WIDTH($signed(P[4151-:32]) / 8)) HWSTRBReg(
				.clk(HCLK),
				.en(HREADY),
				.d(BusByteMaskM[($signed(P[4151-:32]) / 8) - 1:0]),
				.q(HWSTRB)
			);
		end
	endgenerate
	buscachefsm #(
		.BeatCountThreshold(BeatCountThreshold),
		.AHBWLOGBWPL(AHBWLOGBWPL),
		.READ_ONLY_CACHE(READ_ONLY_CACHE),
		.BURST_EN(P[4087])
	) AHBBuscachefsm(
		.HCLK(HCLK),
		.HRESETn(HRESETn),
		.Flush(Flush),
		.BusRW(BusRW),
		.BusAtomic(BusAtomic),
		.Stall(Stall),
		.BusCommitted(BusCommitted),
		.BusStall(BusStall),
		.CaptureEn(CaptureEn),
		.SelBusBeat(SelBusBeat),
		.CacheBusRW(CacheBusRW),
		.BusCMOZero(BusCMOZero),
		.CacheBusAck(CacheBusAck),
		.BeatCount(BeatCount),
		.BeatCountDelayed(BeatCountDelayed),
		.HREADY(HREADY),
		.HTRANS(HTRANS),
		.HWRITE(HWRITE),
		.HBURST(HBURST)
	);
endmodule
module ahbinterface (
	HCLK,
	HRESETn,
	HREADY,
	HTRANS,
	HWRITE,
	HRDATA,
	HWDATA,
	HWSTRB,
	Stall,
	Flush,
	BusRW,
	BusAtomic,
	ByteMask,
	WriteData,
	BusStall,
	BusCommitted,
	FetchBuffer
);
	parameter XLEN = 0;
	parameter [0:0] LSU = 1'b0;
	input wire HCLK;
	input wire HRESETn;
	input wire HREADY;
	output wire [1:0] HTRANS;
	output wire HWRITE;
	input wire [XLEN - 1:0] HRDATA;
	output wire [XLEN - 1:0] HWDATA;
	output wire [(XLEN / 8) - 1:0] HWSTRB;
	input wire Stall;
	input wire Flush;
	input wire [1:0] BusRW;
	input wire BusAtomic;
	input wire [(XLEN / 8) - 1:0] ByteMask;
	input wire [XLEN - 1:0] WriteData;
	output wire BusStall;
	output wire BusCommitted;
	output wire [XLEN - 1:0] FetchBuffer;
	wire CaptureEn;
	flopen #(.WIDTH(XLEN)) fb(
		.clk(HCLK),
		.en(CaptureEn),
		.d(HRDATA),
		.q(FetchBuffer)
	);
	generate
		if (LSU) begin : genblk1
			flop #(.WIDTH(XLEN)) wdreg(
				.clk(HCLK),
				.d(WriteData),
				.q(HWDATA)
			);
			flop #(.WIDTH(XLEN / 8)) HWSTRBReg(
				.clk(HCLK),
				.d(ByteMask),
				.q(HWSTRB)
			);
		end
		else begin : genblk1
			assign HWDATA = 1'sb0;
			assign HWSTRB = 1'sb0;
		end
	endgenerate
	busfsm #(.READ_ONLY(~LSU)) busfsm(
		.HCLK(HCLK),
		.HRESETn(HRESETn),
		.Flush(Flush),
		.BusRW(BusRW),
		.BusAtomic(BusAtomic),
		.BusCommitted(BusCommitted),
		.Stall(Stall),
		.BusStall(BusStall),
		.CaptureEn(CaptureEn),
		.HREADY(HREADY),
		.HTRANS(HTRANS),
		.HWRITE(HWRITE)
	);
endmodule
module buscachefsm (
	HCLK,
	HRESETn,
	Stall,
	Flush,
	BusRW,
	BusAtomic,
	BusCMOZero,
	BusStall,
	BusCommitted,
	CaptureEn,
	CacheBusRW,
	CacheBusAck,
	BeatCount,
	BeatCountDelayed,
	SelBusBeat,
	HREADY,
	HTRANS,
	HWRITE,
	HBURST
);
	reg _sv2v_0;
	parameter BeatCountThreshold = 0;
	parameter AHBWLOGBWPL = 0;
	parameter READ_ONLY_CACHE = 0;
	parameter BURST_EN = 0;
	input wire HCLK;
	input wire HRESETn;
	input wire Stall;
	input wire Flush;
	input wire [1:0] BusRW;
	input wire BusAtomic;
	input wire BusCMOZero;
	output wire BusStall;
	output wire BusCommitted;
	output wire CaptureEn;
	input wire [1:0] CacheBusRW;
	output wire CacheBusAck;
	output wire [AHBWLOGBWPL - 1:0] BeatCount;
	output wire [AHBWLOGBWPL - 1:0] BeatCountDelayed;
	output wire SelBusBeat;
	input wire HREADY;
	output wire [1:0] HTRANS;
	output wire HWRITE;
	output wire [2:0] HBURST;
	reg [2:0] CurrState;
	reg [2:0] NextState;
	wire [AHBWLOGBWPL - 1:0] NextBeatCount;
	wire FinalBeatCount;
	reg [2:0] LocalBurstType;
	wire BeatCntEn;
	wire BeatCntReset;
	wire CacheAccess;
	wire BusWrite;
	assign BusWrite = (CacheBusRW[0] | BusCMOZero) & ~READ_ONLY_CACHE;
	always @(posedge HCLK)
		if (~HRESETn | Flush)
			CurrState <= 3'd0;
		else
			CurrState <= NextState;
	always @(*) begin
		if (_sv2v_0)
			;
		case (CurrState)
			3'd0:
				if (HREADY & |BusRW)
					NextState = 3'd1;
				else if ((HREADY & BusWrite) & ~READ_ONLY_CACHE)
					NextState = 3'd6;
				else if (HREADY & CacheBusRW[1])
					NextState = 3'd5;
				else
					NextState = 3'd0;
			3'd1:
				if ((HREADY & BusAtomic) & ~READ_ONLY_CACHE)
					NextState = 3'd2;
				else if (HREADY & ~BusAtomic)
					NextState = 3'd4;
				else
					NextState = 3'd1;
			3'd2:
				if (HREADY)
					NextState = 3'd3;
				else
					NextState = 3'd2;
			3'd3:
				if (HREADY)
					NextState = 3'd4;
				else
					NextState = 3'd3;
			3'd4:
				if (Stall)
					NextState = 3'd4;
				else
					NextState = 3'd0;
			3'd5:
				if ((HREADY & FinalBeatCount) & CacheBusRW[0])
					NextState = 3'd6;
				else if ((HREADY & FinalBeatCount) & CacheBusRW[1])
					NextState = 3'd5;
				else if ((HREADY & FinalBeatCount) & ~|CacheBusRW)
					NextState = 3'd0;
				else
					NextState = 3'd5;
			3'd6:
				if ((HREADY & FinalBeatCount) & CacheBusRW[0])
					NextState = 3'd6;
				else if ((HREADY & FinalBeatCount) & CacheBusRW[1])
					NextState = 3'd5;
				else if ((HREADY & FinalBeatCount) & BusCMOZero)
					NextState = 3'd4;
				else if ((HREADY & FinalBeatCount) & ~|CacheBusRW)
					NextState = 3'd0;
				else
					NextState = 3'd6;
			default: NextState = 3'd0;
		endcase
	end
	flopenr #(.WIDTH(AHBWLOGBWPL)) BeatCountReg(
		.clk(HCLK),
		.reset(~HRESETn | BeatCntReset),
		.en(BeatCntEn),
		.d(NextBeatCount),
		.q(BeatCount)
	);
	flopenr #(.WIDTH(AHBWLOGBWPL)) BeatCountDelayedReg(
		.clk(HCLK),
		.reset(~HRESETn | BeatCntReset),
		.en(BeatCntEn),
		.d(BeatCount),
		.q(BeatCountDelayed)
	);
	assign NextBeatCount = BeatCount + 1'b1;
	assign FinalBeatCount = BeatCountDelayed == BeatCountThreshold[AHBWLOGBWPL - 1:0];
	assign BeatCntEn = (((((NextState == 3'd6) | (NextState == 3'd5)) & HREADY) & ~Flush) | (((NextState == 3'd0) & |CacheBusRW) & HREADY)) & ~Flush;
	assign BeatCntReset = NextState == 3'd0;
	assign CaptureEn = (((CurrState == 3'd1) & BusRW[1]) & ~Flush) | ((CurrState == 3'd5) & HREADY);
	assign CacheAccess = (CurrState == 3'd5) | (CurrState == 3'd6);
	assign BusStall = ((((((CurrState == 3'd0) & ((|BusRW | (|CacheBusRW)) | BusCMOZero)) | (CurrState == 3'd1)) | (CurrState == 3'd3)) | (CurrState == 3'd2)) | ((CurrState == 3'd5) & ~FinalBeatCount)) | ((CurrState == 3'd6) & ~FinalBeatCount);
	assign BusCommitted = (CurrState != 3'd0) & ~(READ_ONLY_CACHE & (CurrState == 3'd4));
	assign HTRANS = ((((((CurrState == 3'd0) & HREADY) & ((|BusRW | (|CacheBusRW)) | BusCMOZero)) & ~Flush) | (CurrState == 3'd2)) | ((((CacheAccess & FinalBeatCount) & |CacheBusRW) & HREADY) & ~Flush) ? 2'b10 : (CacheAccess & |BeatCount ? (BURST_EN ? 2'b11 : 2'b10) : 2'b00));
	assign HWRITE = ((((BusRW[0] & ~BusAtomic) | (BusWrite & ~Flush)) | ((CurrState == 3'd2) & BusAtomic)) | ((CurrState == 3'd6) & |BeatCount)) & ~READ_ONLY_CACHE;
	assign HBURST = (BURST_EN & ((|CacheBusRW & ~Flush) | (CacheAccess & |BeatCount)) ? LocalBurstType : 3'b000);
	always @(*) begin
		if (_sv2v_0)
			;
		case (BeatCountThreshold)
			0: LocalBurstType = 3'b000;
			3: LocalBurstType = 3'b011;
			7: LocalBurstType = 3'b101;
			15: LocalBurstType = 3'b111;
			default: LocalBurstType = 3'b001;
		endcase
	end
	assign CacheBusAck = ((CacheAccess & HREADY) & FinalBeatCount) & ~BusCMOZero;
	assign SelBusBeat = ((((((CurrState == 3'd0) & (BusRW[0] | BusWrite)) | ((CurrState == 3'd1) & BusRW[0])) | ((CurrState == 3'd3) & BusRW[0])) | ((CurrState == 3'd2) & BusRW[0])) | (CurrState == 3'd6)) | (CurrState == 3'd5);
	initial _sv2v_0 = 0;
endmodule
module busfsm (
	HCLK,
	HRESETn,
	Stall,
	Flush,
	BusRW,
	BusAtomic,
	CaptureEn,
	BusStall,
	BusCommitted,
	HREADY,
	HTRANS,
	HWRITE
);
	reg _sv2v_0;
	parameter [0:0] READ_ONLY = 0;
	input wire HCLK;
	input wire HRESETn;
	input wire Stall;
	input wire Flush;
	input wire [1:0] BusRW;
	input wire BusAtomic;
	output wire CaptureEn;
	output wire BusStall;
	output wire BusCommitted;
	input wire HREADY;
	output wire [1:0] HTRANS;
	output wire HWRITE;
	reg [2:0] CurrState;
	reg [2:0] NextState;
	always @(posedge HCLK)
		if (~HRESETn | Flush)
			CurrState <= 3'd0;
		else
			CurrState <= NextState;
	always @(*) begin
		if (_sv2v_0)
			;
		case (CurrState)
			3'd0:
				if (HREADY & |BusRW)
					NextState = 3'd1;
				else
					NextState = 3'd0;
			3'd1:
				if (HREADY & BusAtomic)
					NextState = 3'd3;
				else if (HREADY & ~BusAtomic)
					NextState = 3'd2;
				else
					NextState = 3'd1;
			3'd3:
				if (HREADY)
					NextState = 3'd4;
				else
					NextState = 3'd3;
			3'd4:
				if (HREADY)
					NextState = 3'd2;
				else
					NextState = 3'd4;
			3'd2:
				if (Stall)
					NextState = 3'd2;
				else
					NextState = 3'd0;
			default: NextState = 3'd0;
		endcase
	end
	assign BusStall = ((((CurrState == 3'd0) & |BusRW) | (CurrState == 3'd4)) | (CurrState == 3'd3)) | (CurrState == 3'd1);
	assign BusCommitted = (CurrState != 3'd0) & ~(READ_ONLY & (CurrState == 3'd2));
	assign HTRANS = (((((CurrState == 3'd0) & HREADY) & |BusRW) & ~Flush) | ((CurrState == 3'd3) & BusAtomic) ? 2'b10 : 2'b00);
	assign HWRITE = (BusRW[0] & ~BusAtomic) | ((CurrState == 3'd3) & BusAtomic);
	assign CaptureEn = CurrState == 3'd1;
	initial _sv2v_0 = 0;
endmodule
module controllerinput (
	HCLK,
	HRESETn,
	Save,
	Restore,
	Disable,
	Request,
	HTRANSIn,
	HWRITEIn,
	HSIZEIn,
	HBURSTIn,
	HADDRIn,
	HREADYOut,
	HTRANSOut,
	HWRITEOut,
	HSIZEOut,
	HBURSTOut,
	HADDROut,
	HREADYIn
);
	parameter PA_BITS = 0;
	parameter SAVE_ENABLED = 1;
	input wire HCLK;
	input wire HRESETn;
	input wire Save;
	input wire Restore;
	input wire Disable;
	output wire Request;
	input wire [1:0] HTRANSIn;
	input wire HWRITEIn;
	input wire [2:0] HSIZEIn;
	input wire [2:0] HBURSTIn;
	input wire [PA_BITS - 1:0] HADDRIn;
	output wire HREADYOut;
	output wire [1:0] HTRANSOut;
	output wire HWRITEOut;
	output wire [2:0] HSIZEOut;
	output wire [2:0] HBURSTOut;
	output wire [PA_BITS - 1:0] HADDROut;
	input wire HREADYIn;
	wire HWRITESave;
	wire [2:0] HSIZESave;
	wire [2:0] HBURSTSave;
	wire [1:0] HTRANSSave;
	wire [PA_BITS - 1:0] HADDRSave;
	generate
		if (SAVE_ENABLED) begin : genblk1
			flopenr #(.WIDTH(9 + PA_BITS)) SaveReg(
				.clk(HCLK),
				.reset(~HRESETn),
				.en(Save),
				.d({HWRITEIn, HSIZEIn, HBURSTIn, HTRANSIn, HADDRIn}),
				.q({HWRITESave, HSIZESave, HBURSTSave, HTRANSSave, HADDRSave})
			);
			mux2 #(.WIDTH(9 + PA_BITS)) RestorMux(
				.d0({HWRITEIn, HSIZEIn, HBURSTIn, HTRANSIn, HADDRIn}),
				.d1({HWRITESave, HSIZESave, HBURSTSave, HTRANSSave, HADDRSave}),
				.s(Restore),
				.y({HWRITEOut, HSIZEOut, HBURSTOut, HTRANSOut, HADDROut})
			);
		end
		else begin : genblk1
			assign HWRITEOut = HWRITEIn;
			assign HSIZEOut = HSIZEIn;
			assign HBURSTOut = HBURSTIn;
			assign HTRANSOut = HTRANSIn;
			assign HADDROut = HADDRIn;
		end
	endgenerate
	assign Request = HTRANSOut != 2'b00;
	assign HREADYOut = HREADYIn & ~Disable;
endmodule
module ebu (
	clk,
	reset,
	IFUHTRANS,
	IFUHSIZE,
	IFUHBURST,
	IFUHADDR,
	IFUHREADY,
	LSUHTRANS,
	LSUHWRITE,
	LSUHSIZE,
	LSUHBURST,
	LSUHADDR,
	LSUHWDATA,
	LSUHWSTRB,
	LSUHREADY,
	HCLK,
	HRESETn,
	HREADY,
	HRESP,
	HADDR,
	HWDATA,
	HWSTRB,
	HWRITE,
	HSIZE,
	HBURST,
	HPROT,
	HTRANS,
	HMASTLOCK
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire [1:0] IFUHTRANS;
	input wire [2:0] IFUHSIZE;
	input wire [2:0] IFUHBURST;
	input wire [$signed(P[1640-:32]) - 1:0] IFUHADDR;
	output wire IFUHREADY;
	input wire [1:0] LSUHTRANS;
	input wire LSUHWRITE;
	input wire [2:0] LSUHSIZE;
	input wire [2:0] LSUHBURST;
	input wire [$signed(P[1640-:32]) - 1:0] LSUHADDR;
	input wire [$signed(P[4216-:32]) - 1:0] LSUHWDATA;
	input wire [($signed(P[4216-:32]) / 8) - 1:0] LSUHWSTRB;
	output wire LSUHREADY;
	output wire HCLK;
	output wire HRESETn;
	input wire HREADY;
	input wire HRESP;
	output wire [$signed(P[1640-:32]) - 1:0] HADDR;
	output wire [$signed(P[4151-:32]) - 1:0] HWDATA;
	output wire [($signed(P[4216-:32]) / 8) - 1:0] HWSTRB;
	output wire HWRITE;
	output wire [2:0] HSIZE;
	output wire [2:0] HBURST;
	output wire [3:0] HPROT;
	output wire [1:0] HTRANS;
	output wire HMASTLOCK;
	wire LSUDisable;
	wire LSUSelect;
	wire IFUSave;
	wire IFURestore;
	wire IFUDisable;
	wire IFUSelect;
	wire [$signed(P[1640-:32]) - 1:0] IFUHADDROut;
	wire [1:0] IFUHTRANSOut;
	wire [2:0] IFUHBURSTOut;
	wire [2:0] IFUHSIZEOut;
	wire IFUHWRITEOut;
	wire [$signed(P[1640-:32]) - 1:0] LSUHADDROut;
	wire [1:0] LSUHTRANSOut;
	wire [2:0] LSUHBURSTOut;
	wire [2:0] LSUHSIZEOut;
	wire LSUHWRITEOut;
	wire IFUReq;
	wire LSUReq;
	assign HCLK = clk;
	assign HRESETn = ~reset;
	controllerinput #(.PA_BITS($signed(P[1640-:32]))) IFUInput(
		.HCLK(HCLK),
		.HRESETn(HRESETn),
		.Save(IFUSave),
		.Restore(IFURestore),
		.Disable(IFUDisable),
		.Request(IFUReq),
		.HWRITEIn(1'b0),
		.HSIZEIn(IFUHSIZE),
		.HBURSTIn(IFUHBURST),
		.HTRANSIn(IFUHTRANS),
		.HADDRIn(IFUHADDR),
		.HWRITEOut(IFUHWRITEOut),
		.HSIZEOut(IFUHSIZEOut),
		.HBURSTOut(IFUHBURSTOut),
		.HREADYOut(IFUHREADY),
		.HTRANSOut(IFUHTRANSOut),
		.HADDROut(IFUHADDROut),
		.HREADYIn(HREADY)
	);
	controllerinput #(
		.PA_BITS($signed(P[1640-:32])),
		.SAVE_ENABLED(0)
	) LSUInput(
		.HCLK(HCLK),
		.HRESETn(HRESETn),
		.Save(1'b0),
		.Restore(1'b0),
		.Disable(LSUDisable),
		.Request(LSUReq),
		.HWRITEIn(LSUHWRITE),
		.HSIZEIn(LSUHSIZE),
		.HBURSTIn(LSUHBURST),
		.HTRANSIn(LSUHTRANS),
		.HADDRIn(LSUHADDR),
		.HREADYOut(LSUHREADY),
		.HWRITEOut(LSUHWRITEOut),
		.HSIZEOut(LSUHSIZEOut),
		.HBURSTOut(LSUHBURSTOut),
		.HTRANSOut(LSUHTRANSOut),
		.HADDROut(LSUHADDROut),
		.HREADYIn(HREADY)
	);
	assign HADDR = (LSUSelect ? LSUHADDROut : (IFUSelect ? IFUHADDROut : {$signed(P[1640-:32]) {1'sb0}}));
	assign HSIZE = (LSUSelect ? LSUHSIZEOut : (IFUSelect ? IFUHSIZEOut : {3 {1'sb0}}));
	assign HBURST = (LSUSelect ? LSUHBURSTOut : (IFUSelect ? IFUHBURSTOut : {3 {1'sb0}}));
	assign HTRANS = (LSUSelect ? LSUHTRANSOut : (IFUSelect ? IFUHTRANSOut : {2 {1'sb0}}));
	assign HWRITE = (LSUSelect ? LSUHWRITEOut : 1'b0);
	assign HPROT = {3'b001, LSUSelect};
	assign HMASTLOCK = 1'b0;
	assign HWDATA = LSUHWDATA;
	assign HWSTRB = LSUHWSTRB;
	ebufsmarb ebufsmarb(
		.HCLK(HCLK),
		.HRESETn(HRESETn),
		.HBURST(HBURST),
		.HREADY(HREADY),
		.LSUReq(LSUReq),
		.IFUReq(IFUReq),
		.IFUSave(IFUSave),
		.IFURestore(IFURestore),
		.IFUDisable(IFUDisable),
		.IFUSelect(IFUSelect),
		.LSUDisable(LSUDisable),
		.LSUSelect(LSUSelect)
	);
endmodule
module ebufsmarb (
	HCLK,
	HRESETn,
	HBURST,
	HREADY,
	LSUReq,
	IFUReq,
	IFUSave,
	IFURestore,
	IFUDisable,
	IFUSelect,
	LSUDisable,
	LSUSelect
);
	reg _sv2v_0;
	input wire HCLK;
	input wire HRESETn;
	input wire [2:0] HBURST;
	input wire HREADY;
	input wire LSUReq;
	input wire IFUReq;
	output wire IFUSave;
	output wire IFURestore;
	output wire IFUDisable;
	output wire IFUSelect;
	output wire LSUDisable;
	output wire LSUSelect;
	wire [1:0] CurrState;
	reg [1:0] NextState;
	wire both;
	wire IFUReqDelay;
	wire FinalBeat;
	wire FinalBeatD;
	wire BeatCntEn;
	wire [3:0] BeatCount;
	wire BeatCntReset;
	reg [3:0] Threshold;
	assign both = LSUReq & IFUReq;
	flopenl_8C148 busreg(
		.clk(HCLK),
		.load(~HRESETn),
		.en(1'b1),
		.d(NextState),
		.val(2'd0),
		.q(CurrState)
	);
	always @(*) begin
		if (_sv2v_0)
			;
		case (CurrState)
			2'd0:
				if (both)
					NextState = 2'd1;
				else
					NextState = 2'd0;
			2'd1:
				if ((HREADY & FinalBeatD) & ~(LSUReq & IFUReq))
					NextState = 2'd0;
				else
					NextState = 2'd1;
			default: NextState = 2'd0;
		endcase
	end
	assign IFUSave = (CurrState == 2'd0) & both;
	assign IFURestore = CurrState == 2'd1;
	assign IFUDisable = CurrState == 2'd1;
	assign IFUSelect = (NextState == 2'd1 ? 1'b0 : IFUReq);
	flopr #(.WIDTH(1)) ifureqreg(
		.clk(HCLK),
		.reset(~HRESETn),
		.d(IFUReq),
		.q(IFUReqDelay)
	);
	assign LSUDisable = (CurrState == 2'd1 ? 1'b0 : IFUReqDelay & ~(HREADY & FinalBeatD));
	assign LSUSelect = (NextState == 2'd1 ? 1'b1 : LSUReq);
	assign BeatCntReset = NextState == 2'd0;
	assign FinalBeat = BeatCount == Threshold;
	assign BeatCntEn = (NextState == 2'd1) & HREADY;
	counter #(.WIDTH(4)) BeatCounter(
		.clk(HCLK),
		.reset((~HRESETn | BeatCntReset) | FinalBeat),
		.en(BeatCntEn),
		.q(BeatCount)
	);
	flopenr #(.WIDTH(1)) FinalBeatReg(
		.clk(HCLK),
		.reset(~HRESETn | BeatCntReset),
		.en(BeatCntEn),
		.d(FinalBeat),
		.q(FinalBeatD)
	);
	always @(*) begin
		if (_sv2v_0)
			;
		if (HBURST[2:1] == 2'b00)
			Threshold = 4'b0000;
		else
			Threshold = ('d2 << HBURST[2:1]) - 'd1;
	end
	initial _sv2v_0 = 0;
endmodule
module fclassify (
	Xs,
	XNaN,
	XSNaN,
	XSubnorm,
	XZero,
	XInf,
	ClassRes
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire Xs;
	input wire XNaN;
	input wire XSNaN;
	input wire XSubnorm;
	input wire XZero;
	input wire XInf;
	output wire [$signed(P[4216-:32]) - 1:0] ClassRes;
	wire PInf;
	wire PZero;
	wire PNorm;
	wire PSubnorm;
	wire NInf;
	wire NZero;
	wire NNorm;
	wire NSubnorm;
	wire XNorm;
	assign XNorm = ~(((XNaN | XInf) | XSubnorm) | XZero);
	assign PInf = ~Xs & XInf;
	assign NInf = Xs & XInf;
	assign PNorm = ~Xs & XNorm;
	assign NNorm = Xs & XNorm;
	assign PSubnorm = ~Xs & XSubnorm;
	assign NSubnorm = Xs & XSubnorm;
	assign PZero = ~Xs & XZero;
	assign NZero = Xs & XZero;
	assign ClassRes = {{$signed(P[4216-:32]) - 10 {1'b0}}, XNaN & ~XSNaN, XSNaN, PInf, PNorm, PSubnorm, PZero, NZero, NSubnorm, NNorm, NInf};
endmodule
module fcmp (
	Fmt,
	OpCtrl,
	Zfa,
	Xs,
	Ys,
	Xe,
	Ye,
	Xm,
	Ym,
	XZero,
	YZero,
	XNaN,
	YNaN,
	XSNaN,
	YSNaN,
	X,
	Y,
	CmpNV,
	CmpFpRes,
	CmpIntRes
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[707-:32]) - 1:0] Fmt;
	input wire [2:0] OpCtrl;
	input wire Zfa;
	input wire Xs;
	input wire Ys;
	input wire [$signed(P[837-:32]) - 1:0] Xe;
	input wire [$signed(P[837-:32]) - 1:0] Ye;
	input wire [$signed(P[805-:32]):0] Xm;
	input wire [$signed(P[805-:32]):0] Ym;
	input wire XZero;
	input wire YZero;
	input wire XNaN;
	input wire YNaN;
	input wire XSNaN;
	input wire YSNaN;
	input wire [$signed(P[901-:32]) - 1:0] X;
	input wire [$signed(P[901-:32]) - 1:0] Y;
	output reg CmpNV;
	output reg [$signed(P[901-:32]) - 1:0] CmpFpRes;
	output wire [$signed(P[4216-:32]) - 1:0] CmpIntRes;
	wire LTabs;
	wire LT;
	wire EQ;
	reg [$signed(P[901-:32]) - 1:0] NaNRes;
	wire BothZero;
	wire EitherNaN;
	wire EitherSNaN;
	assign LTabs = {1'b0, Xe, Xm} < {1'b0, Ye, Ym};
	assign LT = ((Xs & ~Ys) | (((Xs & Ys) & ~LTabs) & ~EQ)) | ((~Xs & ~Ys) & LTabs);
	assign EQ = X == Y;
	assign BothZero = XZero & YZero;
	assign EitherNaN = XNaN | YNaN;
	assign EitherSNaN = XSNaN | YSNaN;
	always @(*) begin
		if (_sv2v_0)
			;
		casez (OpCtrl[2:0])
			3'b110: CmpNV = EitherSNaN;
			3'b101: CmpNV = EitherSNaN;
			3'b010: CmpNV = EitherSNaN;
			3'b0z1:
				if (P[4069])
					CmpNV = (Zfa ? EitherSNaN : EitherNaN);
				else
					CmpNV = EitherNaN;
			3'b100: CmpNV = 1'b0;
			default: CmpNV = 1'bx;
		endcase
	end
	function automatic signed [(($signed(P[1227-:32]) - 2) >= 0 ? $signed(P[1227-:32]) - 1 : 3 - $signed(P[1227-:32])) - 1:0] sv2v_cast_46E5E_signed;
		input reg signed [(($signed(P[1227-:32]) - 2) >= 0 ? $signed(P[1227-:32]) - 1 : 3 - $signed(P[1227-:32])) - 1:0] inp;
		sv2v_cast_46E5E_signed = inp;
	endfunction
	function automatic signed [(($signed(P[1097-:32]) - 2) >= 0 ? $signed(P[1097-:32]) - 1 : 3 - $signed(P[1097-:32])) - 1:0] sv2v_cast_B8EE9_signed;
		input reg signed [(($signed(P[1097-:32]) - 2) >= 0 ? $signed(P[1097-:32]) - 1 : 3 - $signed(P[1097-:32])) - 1:0] inp;
		sv2v_cast_B8EE9_signed = inp;
	endfunction
	function automatic signed [(($signed(P[967-:32]) - 2) >= 0 ? $signed(P[967-:32]) - 1 : 3 - $signed(P[967-:32])) - 1:0] sv2v_cast_67652_signed;
		input reg signed [(($signed(P[967-:32]) - 2) >= 0 ? $signed(P[967-:32]) - 1 : 3 - $signed(P[967-:32])) - 1:0] inp;
		sv2v_cast_67652_signed = inp;
	endfunction
	function automatic signed [(($signed(P[611-:32]) - 2) >= 0 ? $signed(P[611-:32]) - 1 : 3 - $signed(P[611-:32])) - 1:0] sv2v_cast_B7E13_signed;
		input reg signed [(($signed(P[611-:32]) - 2) >= 0 ? $signed(P[611-:32]) - 1 : 3 - $signed(P[611-:32])) - 1:0] inp;
		sv2v_cast_B7E13_signed = inp;
	endfunction
	function automatic signed [(($signed(P[481-:32]) - 2) >= 0 ? $signed(P[481-:32]) - 1 : 3 - $signed(P[481-:32])) - 1:0] sv2v_cast_E1570_signed;
		input reg signed [(($signed(P[481-:32]) - 2) >= 0 ? $signed(P[481-:32]) - 1 : 3 - $signed(P[481-:32])) - 1:0] inp;
		sv2v_cast_E1570_signed = inp;
	endfunction
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk1
			if (P[4184]) begin : genblk1
				wire [$signed(P[901-:32]):1] sv2v_tmp_DA76B;
				assign sv2v_tmp_DA76B = {Xs, {$signed(P[837-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:0]};
				always @(*) NaNRes = sv2v_tmp_DA76B;
			end
			else begin : genblk1
				wire [$signed(P[901-:32]):1] sv2v_tmp_202EF;
				assign sv2v_tmp_202EF = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, {$signed(P[805-:32]) - 1 {1'b0}}};
				always @(*) NaNRes = sv2v_tmp_202EF;
			end
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk1
			if (P[4184]) begin : genblk1
				wire [$signed(P[901-:32]):1] sv2v_tmp_69C34;
				assign sv2v_tmp_69C34 = (Fmt ? {Xs, {$signed(P[837-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:0]} : {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, Xs, {$signed(P[643-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[611-:32])]});
				always @(*) NaNRes = sv2v_tmp_69C34;
			end
			else begin : genblk1
				wire [$signed(P[901-:32]):1] sv2v_tmp_88663;
				assign sv2v_tmp_88663 = (Fmt ? {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, {$signed(P[805-:32]) - 1 {1'b0}}} : {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 1'b0, {$signed(P[643-:32]) {1'b1}}, 1'b1, sv2v_cast_B7E13_signed(0)});
				always @(*) NaNRes = sv2v_tmp_88663;
			end
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					P[773-:2]:
						if (P[4184])
							NaNRes = {Xs, {$signed(P[837-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:0]};
						else
							NaNRes = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, {$signed(P[805-:32]) - 1 {1'b0}}};
					P[579-:2]:
						if (P[4184])
							NaNRes = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, Xs, {$signed(P[643-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[611-:32])]};
						else
							NaNRes = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 1'b0, {$signed(P[643-:32]) {1'b1}}, 1'b1, sv2v_cast_B7E13_signed(0)};
					P[449-:2]:
						if (P[4184])
							NaNRes = {{$signed(P[901-:32]) - $signed(P[545-:32]) {1'b1}}, Xs, {$signed(P[513-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[481-:32])]};
						else
							NaNRes = {{$signed(P[901-:32]) - $signed(P[545-:32]) {1'b1}}, 1'b0, {$signed(P[513-:32]) {1'b1}}, 1'b1, sv2v_cast_E1570_signed(0)};
					default: NaNRes = {$signed(P[901-:32]) {1'bx}};
				endcase
			end
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					2'h3:
						if (P[4184])
							NaNRes = {Xs, {$signed(P[837-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:0]};
						else
							NaNRes = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, {$signed(P[805-:32]) - 1 {1'b0}}};
					2'h1:
						if (P[4184])
							NaNRes = {{$signed(P[901-:32]) - $signed(P[1291-:32]) {1'b1}}, Xs, {$signed(P[1259-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[1227-:32])]};
						else
							NaNRes = {{$signed(P[901-:32]) - $signed(P[1291-:32]) {1'b1}}, 1'b0, {$signed(P[1259-:32]) {1'b1}}, 1'b1, sv2v_cast_46E5E_signed(0)};
					2'h0:
						if (P[4184])
							NaNRes = {{$signed(P[901-:32]) - $signed(P[1161-:32]) {1'b1}}, Xs, {$signed(P[1129-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[1097-:32])]};
						else
							NaNRes = {{$signed(P[901-:32]) - $signed(P[1161-:32]) {1'b1}}, 1'b0, {$signed(P[1129-:32]) {1'b1}}, 1'b1, sv2v_cast_B8EE9_signed(0)};
					2'h2:
						if (P[4184])
							NaNRes = {{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, Xs, {$signed(P[999-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[967-:32])]};
						else
							NaNRes = {{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, 1'b0, {$signed(P[999-:32]) {1'b1}}, 1'b1, sv2v_cast_67652_signed(0)};
				endcase
			end
		end
	endgenerate
	always @(*) begin
		if (_sv2v_0)
			;
		if (OpCtrl[0]) begin
			if (Zfa & P[4069]) begin
				if (XNaN | YNaN)
					CmpFpRes = NaNRes;
				else if (LT)
					CmpFpRes = Y;
				else
					CmpFpRes = X;
			end
			else if (XNaN) begin
				if (YNaN)
					CmpFpRes = NaNRes;
				else
					CmpFpRes = Y;
			end
			else if (YNaN)
				CmpFpRes = X;
			else if (LT)
				CmpFpRes = Y;
			else
				CmpFpRes = X;
		end
		else if (Zfa & P[4069]) begin
			if (XNaN | YNaN)
				CmpFpRes = NaNRes;
			else if (LT)
				CmpFpRes = X;
			else
				CmpFpRes = Y;
		end
		else if (XNaN) begin
			if (YNaN)
				CmpFpRes = NaNRes;
			else
				CmpFpRes = Y;
		end
		else if (YNaN)
			CmpFpRes = X;
		else if (LT)
			CmpFpRes = X;
		else
			CmpFpRes = Y;
	end
	function automatic signed [(($signed(P[4216-:32]) - 2) >= 0 ? $signed(P[4216-:32]) - 1 : 3 - $signed(P[4216-:32])) - 1:0] sv2v_cast_EFBE2_signed;
		input reg signed [(($signed(P[4216-:32]) - 2) >= 0 ? $signed(P[4216-:32]) - 1 : 3 - $signed(P[4216-:32])) - 1:0] inp;
		sv2v_cast_EFBE2_signed = inp;
	endfunction
	assign CmpIntRes = {sv2v_cast_EFBE2_signed(0), (((EQ | BothZero) & OpCtrl[1]) | ((LT & OpCtrl[0]) & ~BothZero)) & ~EitherNaN};
	initial _sv2v_0 = 0;
endmodule
module fctrl (
	clk,
	reset,
	StallE,
	StallM,
	StallW,
	FlushE,
	FlushM,
	FlushW,
	IntDivE,
	FRM_REGW,
	STATUS_FS,
	FDivBusyE,
	InstrD,
	Funct7D,
	OpD,
	Rs2D,
	Funct3D,
	XEnD,
	YEnD,
	ZEnD,
	XEnE,
	YEnE,
	ZEnE,
	FCvtIntE,
	FCvtIntW,
	FrmE,
	FrmM,
	FmtE,
	FmtM,
	OpCtrlE,
	OpCtrlM,
	FpLoadStoreM,
	PostProcSelE,
	PostProcSelM,
	FResSelE,
	FResSelM,
	FResSelW,
	FPUActiveE,
	ZfaE,
	ZfaM,
	ZfaFRoundNXE,
	FRegWriteE,
	FRegWriteM,
	FRegWriteW,
	FWriteIntE,
	FWriteIntM,
	Adr1D,
	Adr2D,
	Adr3D,
	Adr1E,
	Adr2E,
	Adr3E,
	IllegalFPUInstrD,
	FDivStartE,
	IDivStartE
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	input wire IntDivE;
	input wire [2:0] FRM_REGW;
	input wire [1:0] STATUS_FS;
	input wire FDivBusyE;
	input wire [31:0] InstrD;
	input wire [6:0] Funct7D;
	input wire [6:0] OpD;
	input wire [4:0] Rs2D;
	input wire [2:0] Funct3D;
	output wire XEnD;
	output wire YEnD;
	output wire ZEnD;
	output wire XEnE;
	output wire YEnE;
	output wire ZEnE;
	output wire FCvtIntE;
	output wire FCvtIntW;
	output wire [2:0] FrmE;
	output wire [2:0] FrmM;
	output wire [$signed(P[707-:32]) - 1:0] FmtE;
	output wire [$signed(P[707-:32]) - 1:0] FmtM;
	output wire [2:0] OpCtrlE;
	output wire [2:0] OpCtrlM;
	output wire FpLoadStoreM;
	output wire [1:0] PostProcSelE;
	output wire [1:0] PostProcSelM;
	output wire [1:0] FResSelE;
	output wire [1:0] FResSelM;
	output wire [1:0] FResSelW;
	output wire FPUActiveE;
	output wire ZfaE;
	output wire ZfaM;
	output wire ZfaFRoundNXE;
	output wire FRegWriteE;
	output wire FRegWriteM;
	output wire FRegWriteW;
	output wire FWriteIntE;
	output wire FWriteIntM;
	output wire [4:0] Adr1D;
	output wire [4:0] Adr2D;
	output wire [4:0] Adr3D;
	output wire [4:0] Adr1E;
	output wire [4:0] Adr2E;
	output wire [4:0] Adr3E;
	output wire IllegalFPUInstrD;
	output wire FDivStartE;
	output wire IDivStartE;
	reg [13:0] ControlsD;
	wire FRegWriteD;
	wire FDivStartD;
	wire FWriteIntD;
	wire [2:0] OpCtrlD;
	wire [1:0] PostProcSelD;
	wire [1:0] FResSelD;
	wire [2:0] FrmD;
	wire [$signed(P[707-:32]) - 1:0] FmtD;
	wire [1:0] Fmt;
	wire [1:0] Fmt2;
	wire SupportedFmt;
	wire SupportedFmt2;
	wire SupportedRM;
	wire FCvtIntD;
	wire FCvtIntM;
	wire ZfaD;
	wire ZfaFRoundNXD;
	assign Fmt = Funct7D[1:0];
	assign Fmt2 = Rs2D[1:0];
	assign SupportedFmt = (((Fmt == 2'b00) | ((Fmt == 2'b01) & P[1493])) | ((Fmt == 2'b10) & P[4070])) | ((Fmt == 2'b11) & P[1488]);
	assign SupportedFmt2 = (((Fmt2 == 2'b00) | ((Fmt2 == 2'b01) & P[1493])) | ((Fmt2 == 2'b10) & P[4070])) | ((Fmt2 == 2'b11) & P[1488]);
	assign SupportedRM = ~(((Funct3D == 3'b101) | (Funct3D == 3'b110)) | ((Funct3D == 3'b111) & (((FRM_REGW == 3'b101) | (FRM_REGW == 3'b110)) | (FRM_REGW == 3'b111)))) | ((((OpD == 7'b1010011) & (Funct3D == 3'b101)) & (Funct7D[6:2] == 5'b10100)) & P[4069]);
	always @(*) begin
		if (_sv2v_0)
			;
		if (STATUS_FS == 2'b00)
			ControlsD = 14'b00000000001000;
		else if (((OpD != 7'b0000111) & (OpD != 7'b0100111)) & (~SupportedFmt | ~SupportedRM))
			ControlsD = 14'b00000000001000;
		else begin
			ControlsD = 14'b00000000001000;
			case (OpD)
				7'b0000111:
					case (Funct3D)
						3'b010: ControlsD = 14'b1010000xx00000;
						3'b011:
							if (P[1493])
								ControlsD = 14'b1010000xx00000;
						3'b100:
							if (P[1488])
								ControlsD = 14'b1010000xx00000;
						3'b001:
							if (P[4070])
								ControlsD = 14'b1010000xx00000;
					endcase
				7'b0100111:
					case (Funct3D)
						3'b010: ControlsD = 14'b0010000xx00000;
						3'b011:
							if (P[1493])
								ControlsD = 14'b0010000xx00000;
						3'b100:
							if (P[1488])
								ControlsD = 14'b0010000xx00000;
						3'b001:
							if (P[4070])
								ControlsD = 14'b0010000xx00000;
					endcase
				7'b1000011: ControlsD = 14'b10011000000000;
				7'b1000111: ControlsD = 14'b10011000100000;
				7'b1001011: ControlsD = 14'b10011001000000;
				7'b1001111: ControlsD = 14'b10011001100000;
				7'b1010011:
					casez (Funct7D)
						7'b00000zz: ControlsD = 14'b10011011000000;
						7'b00001zz: ControlsD = 14'b10011011100000;
						7'b00010zz: ControlsD = 14'b10011010000000;
						7'b00011zz: ControlsD = 14'b100101xx010000;
						7'b01011zz:
							if (Rs2D == 5'b00000)
								ControlsD = 14'b100101xx110000;
						7'b00100zz:
							case (Funct3D)
								3'b000: ControlsD = 14'b10000000000000;
								3'b001: ControlsD = 14'b10000000100000;
								3'b010: ControlsD = 14'b10000001000000;
							endcase
						7'b00101zz:
							case (Funct3D)
								3'b000: ControlsD = 14'b10000011000000;
								3'b001: ControlsD = 14'b10000010100000;
								3'b010:
									if (P[4069])
										ControlsD = 14'b10000011000010;
								3'b011:
									if (P[4069])
										ControlsD = 14'b10000010100010;
							endcase
						7'b10100zz:
							case (Funct3D)
								3'b000: ControlsD = 14'b01000001100000;
								3'b001: ControlsD = 14'b01000000100000;
								3'b010: ControlsD = 14'b01000001000000;
								3'b100:
									if (P[4069])
										ControlsD = 14'b01000001100010;
								3'b101:
									if (P[4069])
										ControlsD = 14'b01000000100010;
							endcase
						7'b11100zz:
							if ((Funct3D == 3'b001) & (Rs2D == 5'b00000))
								ControlsD = 14'b01100000000000;
							else if ((Funct3D == 3'b000) & (Rs2D == 5'b00000)) begin
								if (((Fmt[1:0] == 2'b00) | (Fmt[1:0] == 2'b10)) | (($signed(P[4216-:32]) == 64) & (Fmt[1:0] == 2'b01)))
									ControlsD = 14'b01110000000000;
							end
							else if (((((P[4069] & ($signed(P[4216-:32]) == 32)) & P[1493]) & (Funct7D[1:0] == 2'b01)) & (Funct3D == 3'b000)) & (Rs2D == 5'b00001))
								ControlsD = 14'b01110000000010;
							else if (((((P[4069] & ($signed(P[4216-:32]) == 64)) & P[1488]) & (Funct7D[1:0] == 2'b11)) & (Funct3D == 3'b000)) & (Rs2D == 5'b00001))
								ControlsD = 14'b01110000000010;
						7'b11110zz:
							if ((Funct3D == 3'b000) & (Rs2D == 5'b00000)) begin
								if (((Fmt[1:0] == 2'b00) | (Fmt[1:0] == 2'b10)) | (($signed(P[4216-:32]) == 64) & (Fmt[1:0] == 2'b01)))
									ControlsD = 14'b10000001100000;
							end
							else if ((P[4069] & (Funct3D == 3'b000)) & (Rs2D == 5'b00001))
								ControlsD = 14'b10000011100010;
						7'b0100000:
							if (((Rs2D[4:2] == 3'b000) & SupportedFmt2) & (Rs2D[1:0] != 2'b00))
								ControlsD = 14'b10010000000000;
							else if ((Rs2D == 5'b00100) & P[4069])
								ControlsD = 14'b10000010000010;
							else if ((Rs2D == 5'b00101) & P[4069])
								ControlsD = 14'b10000010000011;
						7'b0100001:
							if (((Rs2D[4:2] == 3'b000) & SupportedFmt2) & (Rs2D[1:0] != 2'b01))
								ControlsD = 14'b10010000100000;
							else if ((Rs2D == 5'b00100) & P[4069])
								ControlsD = 14'b10000010000010;
							else if ((Rs2D == 5'b00101) & P[4069])
								ControlsD = 14'b10000010000011;
						7'b0100010:
							if (((Rs2D[4:2] == 3'b000) & SupportedFmt2) & (Rs2D[1:0] != 2'b10))
								ControlsD = 14'b10010001000000;
							else if ((Rs2D == 5'b00100) & P[4069])
								ControlsD = 14'b10000010000010;
							else if ((Rs2D == 5'b00101) & P[4069])
								ControlsD = 14'b10000010000011;
						7'b0100011:
							if (((Rs2D[4:2] == 3'b000) & SupportedFmt2) & (Rs2D[1:0] != 2'b11))
								ControlsD = 14'b10010001100000;
							else if ((Rs2D == 5'b00100) & P[4069])
								ControlsD = 14'b10000010000010;
							else if ((Rs2D == 5'b00101) & P[4069])
								ControlsD = 14'b10000010000011;
						7'b1101000:
							case (Rs2D)
								5'b00000: ControlsD = 14'b10010010100000;
								5'b00001: ControlsD = 14'b10010010000000;
								5'b00010:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b10010011100000;
								5'b00011:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b10010011000000;
							endcase
						7'b1100000:
							case (Rs2D)
								5'b00000: ControlsD = 14'b01010000100100;
								5'b00001: ControlsD = 14'b01010000000100;
								5'b00010:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b01010001100100;
								5'b00011:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b01010001000100;
							endcase
						7'b1101001:
							case (Rs2D)
								5'b00000: ControlsD = 14'b10010010100000;
								5'b00001: ControlsD = 14'b10010010000000;
								5'b00010:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b10010011100000;
								5'b00011:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b10010011000000;
							endcase
						7'b1100001:
							case (Rs2D)
								5'b00000: ControlsD = 14'b01010000100100;
								5'b00001: ControlsD = 14'b01010000000100;
								5'b00010:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b01010001100100;
								5'b00011:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b01010001000100;
								5'b01000:
									if ((P[4069] & P[1493]) & (Funct3D == 3'b001))
										ControlsD = 14'b01010000100110;
							endcase
						7'b1101010:
							case (Rs2D)
								5'b00000: ControlsD = 14'b10010010100000;
								5'b00001: ControlsD = 14'b10010010000000;
								5'b00010:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b10010011100000;
								5'b00011:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b10010011000000;
							endcase
						7'b1100010:
							case (Rs2D)
								5'b00000: ControlsD = 14'b01010000100100;
								5'b00001: ControlsD = 14'b01010000000100;
								5'b00010:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b01010001100100;
								5'b00011:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b01010001000100;
							endcase
						7'b1101011:
							case (Rs2D)
								5'b00000: ControlsD = 14'b10010010100000;
								5'b00001: ControlsD = 14'b10010010000000;
								5'b00010:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b10010011100000;
								5'b00011:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b10010011000000;
							endcase
						7'b1100011:
							case (Rs2D)
								5'b00000: ControlsD = 14'b01010000100100;
								5'b00001: ControlsD = 14'b01010000000100;
								5'b00010:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b01010001100100;
								5'b00011:
									if ($signed(P[4216-:32]) == 64)
										ControlsD = 14'b01010001000100;
							endcase
						7'b1011001:
							if (((P[4069] & ($signed(P[4216-:32]) == 32)) & P[1493]) & (Funct3D == 3'b000))
								ControlsD = 14'b10000001100010;
						7'b1011011:
							if (((P[4069] & ($signed(P[4216-:32]) == 64)) & P[1488]) & (Funct3D == 3'b000))
								ControlsD = 14'b10000001100010;
					endcase
			endcase
		end
	end
	assign {FRegWriteD, FWriteIntD, FResSelD, PostProcSelD, OpCtrlD, FDivStartD, IllegalFPUInstrD, FCvtIntD, ZfaD, ZfaFRoundNXD} = ControlsD;
	assign FrmD = (Funct3D == 3'b111 ? FRM_REGW : Funct3D);
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk1
			assign FmtD = 1'b0;
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk1
			wire [1:0] FmtTmp;
			assign FmtTmp = (((Funct7D[6:3] == 4'b0100) & OpD[4]) & ~Rs2D[2] ? Rs2D[1:0] : (~OpD[6] & (&OpD[2:0]) ? {~Funct3D[1], ~(Funct3D[1] ^ Funct3D[0])} : Funct7D[1:0]));
			assign FmtD = P[773-:2] == FmtTmp;
		end
		else if (($signed(P[739-:32]) == 3) | ($signed(P[739-:32]) == 4)) begin : genblk1
			assign FmtD = (((Funct7D[6:3] == 4'b0100) & OpD[4]) & ~Rs2D[2] ? Rs2D[1:0] : Funct7D[1:0]);
		end
	endgenerate
	assign XEnD = ~((((FResSelD == 2'b10) & ~FWriteIntD) | (((FResSelD == 2'b00) & FRegWriteD) & (OpCtrlD == 3'b011))) | (((FResSelD == 2'b01) & (PostProcSelD == 2'b00)) & OpCtrlD[2]));
	assign YEnD = ~(((((FResSelD == 2'b10) & (FWriteIntD | FRegWriteD)) | (((FResSelD == 2'b00) & FRegWriteD) & (OpCtrlD == 3'b011))) | ((FResSelD == 2'b11) & (PostProcSelD == 2'b00))) | ((FResSelD == 2'b01) & ((PostProcSelD == 2'b00) | ((PostProcSelD == 2'b01) & OpCtrlD[0]))));
	assign ZEnD = (PostProcSelD == 2'b10) & (~OpCtrlD[2] | OpCtrlD[1]);
	assign Adr1D = InstrD[19:15];
	assign Adr2D = InstrD[24:20];
	assign Adr3D = InstrD[31:27];
	flopenrc #(.WIDTH(16 + $signed(P[707-:32]))) DECtrlReg3(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d({FRegWriteD, PostProcSelD, FResSelD, FrmD, FmtD, OpCtrlD, FWriteIntD, FCvtIntD, ZfaD, ZfaFRoundNXD, ~IllegalFPUInstrD}),
		.q({FRegWriteE, PostProcSelE, FResSelE, FrmE, FmtE, OpCtrlE, FWriteIntE, FCvtIntE, ZfaE, ZfaFRoundNXE, FPUActiveE})
	);
	flopenrc #(.WIDTH(15)) DEAdrReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d({Adr1D, Adr2D, Adr3D}),
		.q({Adr1E, Adr2E, Adr3E})
	);
	flopenrc #(.WIDTH(1)) DEFDivStartReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE | FDivBusyE),
		.d(FDivStartD),
		.q(FDivStartE)
	);
	flopenrc #(.WIDTH(3)) DEEnReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d({XEnD, YEnD, ZEnD}),
		.q({XEnE, YEnE, ZEnE})
	);
	generate
		if (P[1489] & P[3729]) begin : genblk2
			assign IDivStartE = IntDivE;
		end
		else begin : genblk2
			assign IDivStartE = 1'b0;
		end
	endgenerate
	flopenrc #(.WIDTH(14 + $signed(P[707-:32]))) EMCtrlReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d({FRegWriteE, FResSelE, PostProcSelE, FrmE, FmtE, OpCtrlE, FWriteIntE, FCvtIntE, ZfaE}),
		.q({FRegWriteM, FResSelM, PostProcSelM, FrmM, FmtM, OpCtrlM, FWriteIntM, FCvtIntM, ZfaM})
	);
	assign FpLoadStoreM = FResSelM[1];
	flopenrc #(.WIDTH(4)) MWCtrlReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d({FRegWriteM, FResSelM, FCvtIntM}),
		.q({FRegWriteW, FResSelW, FCvtIntW})
	);
	initial _sv2v_0 = 0;
endmodule
module fcvt (
	Xs,
	Xe,
	Xm,
	Int,
	OpCtrl,
	ToInt,
	XZero,
	Fmt,
	Ce,
	ShiftAmt,
	ResSubnormUf,
	Cs,
	IntZero,
	LzcIn
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire Xs;
	input wire [$signed(P[837-:32]) - 1:0] Xe;
	input wire [$signed(P[805-:32]):0] Xm;
	input wire [$signed(P[4216-:32]) - 1:0] Int;
	input wire [2:0] OpCtrl;
	input wire ToInt;
	input wire XZero;
	input wire [$signed(P[707-:32]) - 1:0] Fmt;
	output wire [$signed(P[837-:32]):0] Ce;
	output reg [$signed(P[351-:32]) - 1:0] ShiftAmt;
	output wire ResSubnormUf;
	output reg Cs;
	output wire IntZero;
	output wire [$signed(P[415-:32]) - 1:0] LzcIn;
	wire [$signed(P[707-:32]) - 1:0] OutFmt;
	wire [$signed(P[4216-:32]) - 1:0] PosInt;
	wire [$signed(P[4216-:32]) - 1:0] TrimInt;
	wire [$signed(P[837-:32]) - 2:0] NewBias;
	wire [$signed(P[837-:32]) - 1:0] OldExp;
	wire Signed;
	wire Int64;
	wire IntToFp;
	wire [$signed(P[415-:32]):0] LzcInFull;
	wire [$signed(P[351-:32]) - 1:0] LeadingZeros;
	assign Signed = OpCtrl[0];
	assign Int64 = OpCtrl[1];
	assign IntToFp = OpCtrl[2];
	generate
		if ($signed(P[739-:32]) == 2) begin : genblk1
			assign OutFmt = (IntToFp ? Fmt : OpCtrl[1:0] == P[773-:2]);
		end
		else if (($signed(P[739-:32]) == 3) | ($signed(P[739-:32]) == 4)) begin : genblk1
			assign OutFmt = (IntToFp ? Fmt : OpCtrl[1:0]);
		end
	endgenerate
	assign PosInt = (Cs ? -Int : Int);
	assign TrimInt = {{$signed(P[4216-:32]) - 32 {Int64}}, {32 {1'b1}}} & PosInt;
	assign IntZero = ~|TrimInt;
	assign LzcInFull = (IntToFp ? {TrimInt, {($signed(P[415-:32]) - $signed(P[4216-:32])) + 1 {1'b0}}} : {Xm, {$signed(P[415-:32]) - $signed(P[805-:32]) {1'b0}}});
	assign LzcIn = LzcInFull[$signed(P[415-:32]) - 1:0];
	lzc #(.WIDTH($signed(P[415-:32]) + 1)) lzc(
		.num(LzcInFull),
		.ZeroCnt(LeadingZeros)
	);
	function automatic signed [(($signed(P[837-:32]) - 2) >= 0 ? $signed(P[837-:32]) - 1 : 3 - $signed(P[837-:32])) - 1:0] sv2v_cast_6B72C_signed;
		input reg signed [(($signed(P[837-:32]) - 2) >= 0 ? $signed(P[837-:32]) - 1 : 3 - $signed(P[837-:32])) - 1:0] inp;
		sv2v_cast_6B72C_signed = inp;
	endfunction
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk2
			assign NewBias = (ToInt ? sv2v_cast_6B72C_signed(1) : sv2v_cast_6B72C_signed($signed(P[771-:32])));
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk2
			reg [$signed(P[837-:32]) - 2:0] NewBiasToFp;
			wire [(($signed(P[837-:32]) - 2) >= 0 ? $signed(P[837-:32]) - 1 : 3 - $signed(P[837-:32])):1] sv2v_tmp_A20ED;
			assign sv2v_tmp_A20ED = (OutFmt ? sv2v_cast_6B72C_signed($signed(P[771-:32])) : sv2v_cast_6B72C_signed($signed(P[577-:32])));
			always @(*) NewBiasToFp = sv2v_tmp_A20ED;
			assign NewBias = (ToInt ? sv2v_cast_6B72C_signed(1) : NewBiasToFp);
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk2
			reg [$signed(P[837-:32]) - 2:0] NewBiasToFp;
			always @(*) begin
				if (_sv2v_0)
					;
				case (OutFmt)
					P[773-:2]: NewBiasToFp = sv2v_cast_6B72C_signed($signed(P[771-:32]));
					P[579-:2]: NewBiasToFp = sv2v_cast_6B72C_signed($signed(P[577-:32]));
					P[449-:2]: NewBiasToFp = sv2v_cast_6B72C_signed($signed(P[447-:32]));
					default: NewBiasToFp = {$signed(P[837-:32]) - 1 {1'bx}};
				endcase
			end
			assign NewBias = (ToInt ? sv2v_cast_6B72C_signed(1) : NewBiasToFp);
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk2
			reg [$signed(P[837-:32]) - 2:0] NewBiasToFp;
			always @(*) begin
				if (_sv2v_0)
					;
				case (OutFmt)
					2'h3: NewBiasToFp = sv2v_cast_6B72C_signed($signed(P[1325-:32]));
					2'h1: NewBiasToFp = sv2v_cast_6B72C_signed($signed(P[1195-:32]));
					2'h0: NewBiasToFp = sv2v_cast_6B72C_signed($signed(P[1065-:32]));
					2'h2: NewBiasToFp = sv2v_cast_6B72C_signed($signed(P[935-:32]));
				endcase
			end
			assign NewBias = (ToInt ? sv2v_cast_6B72C_signed(1) : NewBiasToFp);
		end
	endgenerate
	function automatic signed [$signed(P[837-:32]) - 1:0] sv2v_cast_AF3D4_signed;
		input reg signed [$signed(P[837-:32]) - 1:0] inp;
		sv2v_cast_AF3D4_signed = inp;
	endfunction
	assign OldExp = (IntToFp ? sv2v_cast_AF3D4_signed($signed(P[771-:32])) + sv2v_cast_AF3D4_signed($signed(P[4216-:32]) - 1) : Xe);
	function automatic signed [(($signed(P[837-:32]) + 0) >= 0 ? $signed(P[837-:32]) + 1 : 1 - ($signed(P[837-:32]) + 0)) - 1:0] sv2v_cast_97D7C_signed;
		input reg signed [(($signed(P[837-:32]) + 0) >= 0 ? $signed(P[837-:32]) + 1 : 1 - ($signed(P[837-:32]) + 0)) - 1:0] inp;
		sv2v_cast_97D7C_signed = inp;
	endfunction
	assign Ce = (({1'b0, OldExp} - sv2v_cast_97D7C_signed($signed(P[771-:32]))) - {{($signed(P[837-:32]) - $signed(P[351-:32])) + 1 {1'b0}}, LeadingZeros}) + {2'b00, NewBias};
	assign ResSubnormUf = ((~|Ce | Ce[$signed(P[837-:32])]) & ~XZero) & ~IntToFp;
	function automatic signed [$signed(P[351-:32]) - 1:0] sv2v_cast_AB482_signed;
		input reg signed [$signed(P[351-:32]) - 1:0] inp;
		sv2v_cast_AB482_signed = inp;
	endfunction
	always @(*) begin
		if (_sv2v_0)
			;
		if (ToInt)
			ShiftAmt = Ce[$signed(P[351-:32]) - 1:0] & {$signed(P[351-:32]) {~Ce[$signed(P[837-:32])]}};
		else if (ResSubnormUf)
			ShiftAmt = sv2v_cast_AB482_signed($signed(P[805-:32]) - 1) + Ce[$signed(P[351-:32]) - 1:0];
		else
			ShiftAmt = LeadingZeros;
	end
	always @(*) begin
		if (_sv2v_0)
			;
		if (IntToFp) begin
			if (Int64)
				Cs = Int[$signed(P[4216-:32]) - 1] & Signed;
			else
				Cs = Int[31] & Signed;
		end
		else
			Cs = Xs;
	end
	initial _sv2v_0 = 0;
endmodule
module fhazard (
	Adr1D,
	Adr2D,
	Adr3D,
	Adr1E,
	Adr2E,
	Adr3E,
	FRegWriteE,
	FRegWriteM,
	FRegWriteW,
	RdE,
	RdM,
	RdW,
	FResSelM,
	XEnD,
	YEnD,
	ZEnD,
	FPUStallD,
	ForwardXE,
	ForwardYE,
	ForwardZE
);
	reg _sv2v_0;
	input wire [4:0] Adr1D;
	input wire [4:0] Adr2D;
	input wire [4:0] Adr3D;
	input wire [4:0] Adr1E;
	input wire [4:0] Adr2E;
	input wire [4:0] Adr3E;
	input wire FRegWriteE;
	input wire FRegWriteM;
	input wire FRegWriteW;
	input wire [4:0] RdE;
	input wire [4:0] RdM;
	input wire [4:0] RdW;
	input wire [1:0] FResSelM;
	input wire XEnD;
	input wire YEnD;
	input wire ZEnD;
	output wire FPUStallD;
	output reg [1:0] ForwardXE;
	output reg [1:0] ForwardYE;
	output reg [1:0] ForwardZE;
	wire MatchDE;
	assign MatchDE = (((Adr1D == RdE) & XEnD) | ((Adr2D == RdE) & YEnD)) | ((Adr3D == RdE) & ZEnD);
	assign FPUStallD = MatchDE & FRegWriteE;
	always @(*) begin
		if (_sv2v_0)
			;
		ForwardXE = 2'b00;
		ForwardYE = 2'b00;
		ForwardZE = 2'b00;
		if ((Adr1E == RdM) & FRegWriteM) begin
			if (FResSelM == 2'b00)
				ForwardXE = 2'b10;
		end
		else if ((Adr1E == RdW) & FRegWriteW)
			ForwardXE = 2'b01;
		if ((Adr2E == RdM) & FRegWriteM) begin
			if (FResSelM == 2'b00)
				ForwardYE = 2'b10;
		end
		else if ((Adr2E == RdW) & FRegWriteW)
			ForwardYE = 2'b01;
		if ((Adr3E == RdM) & FRegWriteM) begin
			if (FResSelM == 2'b00)
				ForwardZE = 2'b10;
		end
		else if ((Adr3E == RdW) & FRegWriteW)
			ForwardZE = 2'b01;
	end
	initial _sv2v_0 = 0;
endmodule
module fli (
	Rs1,
	Fmt,
	Imm
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [4:0] Rs1;
	input wire [1:0] Fmt;
	output wire [$signed(P[901-:32]) - 1:0] Imm;
	wire [$signed(P[901-:32]) - 1:0] HImmBox;
	wire [$signed(P[901-:32]) - 1:0] SImmBox;
	wire [$signed(P[901-:32]) - 1:0] DImmBox;
	wire [$signed(P[901-:32]) - 1:0] QImmBox;
	generate
		if (P[4070]) begin : genblk1
			reg [15:0] HImm;
			always @(*) begin
				if (_sv2v_0)
					;
				case (Rs1)
					0: HImm = 16'hbc00;
					1: HImm = 16'h0400;
					2: HImm = 16'h0100;
					3: HImm = 16'h0200;
					4: HImm = 16'h1c00;
					5: HImm = 16'h2000;
					6: HImm = 16'h2c00;
					7: HImm = 16'h3000;
					8: HImm = 16'h3400;
					9: HImm = 16'h3500;
					10: HImm = 16'h3600;
					11: HImm = 16'h3700;
					12: HImm = 16'h3800;
					13: HImm = 16'h3900;
					14: HImm = 16'h3a00;
					15: HImm = 16'h3b00;
					16: HImm = 16'h3c00;
					17: HImm = 16'h3d00;
					18: HImm = 16'h3e00;
					19: HImm = 16'h3f00;
					20: HImm = 16'h4000;
					21: HImm = 16'h4100;
					22: HImm = 16'h4200;
					23: HImm = 16'h4400;
					24: HImm = 16'h4800;
					25: HImm = 16'h4c00;
					26: HImm = 16'h5800;
					27: HImm = 16'h5c00;
					28: HImm = 16'h7800;
					29: HImm = 16'h7c00;
					30: HImm = 16'h7c00;
					31: HImm = 16'h7e00;
				endcase
			end
			assign HImmBox = {{$signed(P[901-:32]) - 16 {1'b1}}, HImm};
		end
		else begin : genblk1
			assign HImmBox = 1'sb0;
		end
	endgenerate
	reg [31:0] SImm;
	always @(*) begin
		if (_sv2v_0)
			;
		case (Rs1)
			0: SImm = 32'hbf800000;
			1: SImm = 32'h00800000;
			2: SImm = 32'h37800000;
			3: SImm = 32'h38000000;
			4: SImm = 32'h3b800000;
			5: SImm = 32'h3c000000;
			6: SImm = 32'h3d800000;
			7: SImm = 32'h3e000000;
			8: SImm = 32'h3e800000;
			9: SImm = 32'h3ea00000;
			10: SImm = 32'h3ec00000;
			11: SImm = 32'h3ee00000;
			12: SImm = 32'h3f000000;
			13: SImm = 32'h3f200000;
			14: SImm = 32'h3f400000;
			15: SImm = 32'h3f600000;
			16: SImm = 32'h3f800000;
			17: SImm = 32'h3fa00000;
			18: SImm = 32'h3fc00000;
			19: SImm = 32'h3fe00000;
			20: SImm = 32'h40000000;
			21: SImm = 32'h40200000;
			22: SImm = 32'h40400000;
			23: SImm = 32'h40800000;
			24: SImm = 32'h41000000;
			25: SImm = 32'h41800000;
			26: SImm = 32'h43000000;
			27: SImm = 32'h43800000;
			28: SImm = 32'h47000000;
			29: SImm = 32'h47800000;
			30: SImm = 32'h7f800000;
			31: SImm = 32'h7fc00000;
		endcase
	end
	assign SImmBox = {{$signed(P[901-:32]) - 32 {1'b1}}, SImm};
	generate
		if (P[1493]) begin : genblk2
			reg [63:0] DImm;
			always @(*) begin
				if (_sv2v_0)
					;
				case (Rs1)
					0: DImm = 64'hbff0000000000000;
					1: DImm = 64'h0010000000000000;
					2: DImm = 64'h3ef0000000000000;
					3: DImm = 64'h3f00000000000000;
					4: DImm = 64'h3f70000000000000;
					5: DImm = 64'h3f80000000000000;
					6: DImm = 64'h3fb0000000000000;
					7: DImm = 64'h3fc0000000000000;
					8: DImm = 64'h3fd0000000000000;
					9: DImm = 64'h3fd4000000000000;
					10: DImm = 64'h3fd8000000000000;
					11: DImm = 64'h3fdc000000000000;
					12: DImm = 64'h3fe0000000000000;
					13: DImm = 64'h3fe4000000000000;
					14: DImm = 64'h3fe8000000000000;
					15: DImm = 64'h3fec000000000000;
					16: DImm = 64'h3ff0000000000000;
					17: DImm = 64'h3ff4000000000000;
					18: DImm = 64'h3ff8000000000000;
					19: DImm = 64'h3ffc000000000000;
					20: DImm = 64'h4000000000000000;
					21: DImm = 64'h4004000000000000;
					22: DImm = 64'h4008000000000000;
					23: DImm = 64'h4010000000000000;
					24: DImm = 64'h4020000000000000;
					25: DImm = 64'h4030000000000000;
					26: DImm = 64'h4060000000000000;
					27: DImm = 64'h4070000000000000;
					28: DImm = 64'h40e0000000000000;
					29: DImm = 64'h40f0000000000000;
					30: DImm = 64'h7ff0000000000000;
					31: DImm = 64'h7ff8000000000000;
				endcase
			end
			assign DImmBox = {{$signed(P[901-:32]) - 64 {1'b1}}, DImm};
		end
		else begin : genblk2
			assign DImmBox = 1'sb0;
		end
		if (P[1488]) begin : genblk3
			reg [127:0] QImm;
			always @(*) begin
				if (_sv2v_0)
					;
				case (Rs1)
					0: QImm = 128'hbfff0000000000000000000000000000;
					1: QImm = 128'h00010000000000000000000000000000;
					2: QImm = 128'h3fef0000000000000000000000000000;
					3: QImm = 128'h3ff00000000000000000000000000000;
					4: QImm = 128'h3ff70000000000000000000000000000;
					5: QImm = 128'h3ff80000000000000000000000000000;
					6: QImm = 128'h3ffb0000000000000000000000000000;
					7: QImm = 128'h3ffc0000000000000000000000000000;
					8: QImm = 128'h3ffd0000000000000000000000000000;
					9: QImm = 128'h3ffd4000000000000000000000000000;
					10: QImm = 128'h3ffd8000000000000000000000000000;
					11: QImm = 128'h3ffdc000000000000000000000000000;
					12: QImm = 128'h3ffe0000000000000000000000000000;
					13: QImm = 128'h3ffe4000000000000000000000000000;
					14: QImm = 128'h3ffe8000000000000000000000000000;
					15: QImm = 128'h3ffec000000000000000000000000000;
					16: QImm = 128'h3fff0000000000000000000000000000;
					17: QImm = 128'h3fff4000000000000000000000000000;
					18: QImm = 128'h3fff8000000000000000000000000000;
					19: QImm = 128'h3fffc000000000000000000000000000;
					20: QImm = 128'h40000000000000000000000000000000;
					21: QImm = 128'h40004000000000000000000000000000;
					22: QImm = 128'h40008000000000000000000000000000;
					23: QImm = 128'h40010000000000000000000000000000;
					24: QImm = 128'h40020000000000000000000000000000;
					25: QImm = 128'h40030000000000000000000000000000;
					26: QImm = 128'h40060000000000000000000000000000;
					27: QImm = 128'h40070000000000000000000000000000;
					28: QImm = 128'h400e0000000000000000000000000000;
					29: QImm = 128'h400f0000000000000000000000000000;
					30: QImm = 128'h7fff0000000000000000000000000000;
					31: QImm = 128'h7fff8000000000000000000000000000;
				endcase
			end
			assign QImmBox = QImm;
		end
		else begin : genblk3
			assign QImmBox = 1'sb0;
		end
	endgenerate
	mux4 #(.WIDTH($signed(P[901-:32]))) flimux(
		.d0(SImmBox),
		.d1(DImmBox),
		.d2(HImmBox),
		.d3(QImmBox),
		.s(Fmt),
		.y(Imm)
	);
	initial _sv2v_0 = 0;
endmodule
module fmtparams (
	Fmt,
	Bias,
	Nf
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[707-:32]) - 1:0] Fmt;
	output reg [$signed(P[837-:32]) - 2:0] Bias;
	output reg [$signed(P[869-:32]) - 1:0] Nf;
	function automatic signed [(($signed(P[837-:32]) - 2) >= 0 ? $signed(P[837-:32]) - 1 : 3 - $signed(P[837-:32])) - 1:0] sv2v_cast_6B72C_signed;
		input reg signed [(($signed(P[837-:32]) - 2) >= 0 ? $signed(P[837-:32]) - 1 : 3 - $signed(P[837-:32])) - 1:0] inp;
		sv2v_cast_6B72C_signed = inp;
	endfunction
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk1
			wire [(($signed(P[837-:32]) - 2) >= 0 ? $signed(P[837-:32]) - 1 : 3 - $signed(P[837-:32])):1] sv2v_tmp_AFE39;
			assign sv2v_tmp_AFE39 = sv2v_cast_6B72C_signed($signed(P[771-:32]));
			always @(*) Bias = sv2v_tmp_AFE39;
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk1
			wire [(($signed(P[837-:32]) - 2) >= 0 ? $signed(P[837-:32]) - 1 : 3 - $signed(P[837-:32])):1] sv2v_tmp_90134;
			assign sv2v_tmp_90134 = (Fmt ? sv2v_cast_6B72C_signed($signed(P[771-:32])) : sv2v_cast_6B72C_signed($signed(P[577-:32])));
			always @(*) Bias = sv2v_tmp_90134;
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					P[773-:2]: Bias = sv2v_cast_6B72C_signed($signed(P[771-:32]));
					P[579-:2]: Bias = sv2v_cast_6B72C_signed($signed(P[577-:32]));
					P[449-:2]: Bias = sv2v_cast_6B72C_signed($signed(P[447-:32]));
					default: Bias = 1'sbx;
				endcase
			end
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					2'h3: Bias = sv2v_cast_6B72C_signed($signed(P[1325-:32]));
					2'h1: Bias = sv2v_cast_6B72C_signed($signed(P[1195-:32]));
					2'h0: Bias = sv2v_cast_6B72C_signed($signed(P[1065-:32]));
					2'h2: Bias = sv2v_cast_6B72C_signed($signed(P[935-:32]));
				endcase
			end
		end
		if ($signed(P[739-:32]) == 1) begin : genblk2
			wire [$signed(P[869-:32]):1] sv2v_tmp_E110F;
			assign sv2v_tmp_E110F = $signed(P[805-:32]);
			always @(*) Nf = sv2v_tmp_E110F;
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk2
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					1'b0: Nf = $signed(P[611-:32]);
					1'b1: Nf = $signed(P[805-:32]);
				endcase
			end
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk2
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					P[773-:2]: Nf = $signed(P[805-:32]);
					P[579-:2]: Nf = $signed(P[611-:32]);
					P[449-:2]: Nf = $signed(P[481-:32]);
					default: Nf = 1'sbx;
				endcase
			end
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk2
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					P[1033-:2]: Nf = $signed(P[1097-:32]);
					P[1163-:2]: Nf = $signed(P[1227-:32]);
					P[903-:2]: Nf = $signed(P[967-:32]);
					P[1293-:2]: Nf = $signed(P[1357-:32]);
				endcase
			end
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module fpu (
	clk,
	reset,
	StallE,
	StallM,
	StallW,
	FlushE,
	FlushM,
	FlushW,
	FPUStallD,
	FDivBusyE,
	STATUS_FS,
	FRM_REGW,
	InstrD,
	Funct3E,
	IntDivE,
	W64E,
	ForwardedSrcAE,
	ForwardedSrcBE,
	RdE,
	FWriteIntE,
	FCvtIntE,
	Funct3M,
	RdM,
	FRegWriteM,
	FpLoadStoreM,
	FWriteDataM,
	FIntResM,
	IllegalFPUInstrD,
	SetFflagsM,
	RdW,
	ReadDataW,
	FCvtIntResW,
	FCvtIntW,
	FIntDivResultW
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	output wire FPUStallD;
	output wire FDivBusyE;
	input wire [1:0] STATUS_FS;
	input wire [2:0] FRM_REGW;
	input wire [31:0] InstrD;
	input wire [2:0] Funct3E;
	input wire IntDivE;
	input wire W64E;
	input wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcAE;
	input wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcBE;
	input wire [4:0] RdE;
	output wire FWriteIntE;
	output wire FCvtIntE;
	input wire [2:0] Funct3M;
	input wire [4:0] RdM;
	output wire FRegWriteM;
	output wire FpLoadStoreM;
	output wire [$signed(P[901-:32]) - 1:0] FWriteDataM;
	output wire [$signed(P[4216-:32]) - 1:0] FIntResM;
	output wire IllegalFPUInstrD;
	output wire [4:0] SetFflagsM;
	input wire [4:0] RdW;
	input wire [$signed(P[901-:32]) - 1:0] ReadDataW;
	output wire [$signed(P[4216-:32]) - 1:0] FCvtIntResW;
	output wire FCvtIntW;
	output wire [$signed(P[4216-:32]) - 1:0] FIntDivResultW;
	wire FRegWriteW;
	wire [2:0] FrmE;
	wire [2:0] FrmM;
	wire [$signed(P[707-:32]) - 1:0] FmtE;
	wire [$signed(P[707-:32]) - 1:0] FmtM;
	wire FDivStartE;
	wire IDivStartE;
	wire FWriteIntM;
	wire [1:0] ForwardXE;
	wire [1:0] ForwardYE;
	wire [1:0] ForwardZE;
	wire [2:0] OpCtrlE;
	wire [2:0] OpCtrlM;
	wire [1:0] FResSelE;
	wire [1:0] FResSelM;
	wire [1:0] FResSelW;
	wire [1:0] PostProcSelE;
	wire [1:0] PostProcSelM;
	wire [4:0] Adr1D;
	wire [4:0] Adr2D;
	wire [4:0] Adr3D;
	wire [4:0] Adr1E;
	wire [4:0] Adr2E;
	wire [4:0] Adr3E;
	wire XEnD;
	wire YEnD;
	wire ZEnD;
	wire XEnE;
	wire YEnE;
	wire ZEnE;
	wire FRegWriteE;
	wire FPUActiveE;
	wire ZfaE;
	wire ZfaM;
	wire ZfaFRoundNXE;
	wire [$signed(P[901-:32]) - 1:0] FRD1D;
	wire [$signed(P[901-:32]) - 1:0] FRD2D;
	wire [$signed(P[901-:32]) - 1:0] FRD3D;
	wire [$signed(P[901-:32]) - 1:0] FRD1E;
	wire [$signed(P[901-:32]) - 1:0] FRD2E;
	wire [$signed(P[901-:32]) - 1:0] FRD3E;
	wire [$signed(P[901-:32]) - 1:0] XE;
	wire [$signed(P[4216-:32]) - 1:0] IntSrcXE;
	wire [$signed(P[901-:32]) - 1:0] PreYE;
	wire [$signed(P[901-:32]) - 1:0] YE;
	wire [$signed(P[901-:32]) - 1:0] PreZE;
	wire [$signed(P[901-:32]) - 1:0] ZE;
	wire XsE;
	wire YsE;
	wire ZsE;
	wire XsM;
	wire YsM;
	wire [$signed(P[837-:32]) - 1:0] XeE;
	wire [$signed(P[837-:32]) - 1:0] YeE;
	wire [$signed(P[837-:32]) - 1:0] ZeE;
	wire [$signed(P[837-:32]) - 1:0] ZeM;
	wire [$signed(P[805-:32]):0] XmE;
	wire [$signed(P[805-:32]):0] YmE;
	wire [$signed(P[805-:32]):0] ZmE;
	wire [$signed(P[805-:32]):0] XmM;
	wire [$signed(P[805-:32]):0] YmM;
	wire [$signed(P[805-:32]):0] ZmM;
	wire XNaNE;
	wire YNaNE;
	wire ZNaNE;
	wire XNaNM;
	wire YNaNM;
	wire ZNaNM;
	wire XSNaNE;
	wire YSNaNE;
	wire ZSNaNE;
	wire XSNaNM;
	wire YSNaNM;
	wire ZSNaNM;
	wire XSubnormE;
	wire XZeroE;
	wire YZeroE;
	wire ZZeroE;
	wire XZeroM;
	wire YZeroM;
	wire XInfE;
	wire YInfE;
	wire ZInfE;
	wire XInfM;
	wire YInfM;
	wire ZInfM;
	wire XExpMaxE;
	wire [$signed(P[901-:32]) - 1:0] XPostBoxE;
	wire [$signed(P[837-:32]) - 2:0] BiasE;
	wire [$signed(P[869-:32]) - 1:0] NfE;
	wire FmaAddSubE;
	wire [1:0] FmaZSelE;
	wire [$signed(P[255-:32]) - 1:0] SmE;
	wire [$signed(P[255-:32]) - 1:0] SmM;
	wire FmaAStickyE;
	wire FmaAStickyM;
	wire [$signed(P[837-:32]) + 1:0] SeE;
	wire [$signed(P[837-:32]) + 1:0] SeM;
	wire InvAE;
	wire InvAM;
	wire AsE;
	wire AsM;
	wire PsE;
	wire PsM;
	wire SsE;
	wire SsM;
	wire [$clog2($signed(P[255-:32]) + 1) - 1:0] SCntE;
	wire [$clog2($signed(P[255-:32]) + 1) - 1:0] SCntM;
	wire [$signed(P[837-:32]):0] CeE;
	wire [$signed(P[837-:32]):0] CeM;
	wire [$signed(P[351-:32]) - 1:0] CvtShiftAmtE;
	wire [$signed(P[351-:32]) - 1:0] CvtShiftAmtM;
	wire CvtResSubnormUfE;
	wire CvtResSubnormUfM;
	wire CsE;
	wire CsM;
	wire IntZeroE;
	wire IntZeroM;
	wire [$signed(P[415-:32]) - 1:0] CvtLzcInE;
	wire [$signed(P[415-:32]) - 1:0] CvtLzcInM;
	wire [$signed(P[4216-:32]) - 1:0] FCvtIntResM;
	wire [$signed(P[95-:32]):0] UmM;
	wire [$signed(P[837-:32]) + 1:0] UeM;
	wire DivStickyM;
	wire FDivDoneE;
	wire IFDivStartE;
	wire [$signed(P[4216-:32]) - 1:0] FIntDivResultM;
	wire [$signed(P[4216-:32]) - 1:0] ClassResE;
	wire [$signed(P[901-:32]) - 1:0] CmpFpResE;
	wire [$signed(P[4216-:32]) - 1:0] CmpIntResE;
	wire CmpNVE;
	wire [$signed(P[901-:32]) - 1:0] SgnResE;
	wire [$signed(P[4216-:32]) - 1:0] FIntResE;
	wire [$signed(P[901-:32]) - 1:0] PostProcResM;
	wire [4:0] PostProcFlgM;
	wire PreNVE;
	wire PreNVM;
	wire PreNXE;
	wire PreNXM;
	wire [$signed(P[901-:32]) - 1:0] FpResM;
	wire [$signed(P[901-:32]) - 1:0] FpResW;
	wire [$signed(P[901-:32]) - 1:0] PreFpResE;
	wire [$signed(P[901-:32]) - 1:0] PreFpResM;
	wire [$signed(P[901-:32]) - 1:0] FResultW;
	wire [$signed(P[901-:32]) - 1:0] PreIntSrcE;
	wire [$signed(P[901-:32]) - 1:0] IntSrcE;
	wire [$signed(P[901-:32]) - 1:0] BoxedZeroE;
	wire [$signed(P[901-:32]) - 1:0] BoxedOneE;
	wire StallUnpackedM;
	wire [$signed(P[901-:32]) - 1:0] SgnExtXE;
	wire mvsgn;
	wire [$signed(P[901-:32]) - 1:0] ZfaResE;
	wire FRoundNVE;
	wire FRoundNXE;
	fctrl #(.P(P)) fctrl(
		.Funct7D(InstrD[31:25]),
		.OpD(InstrD[6:0]),
		.Rs2D(InstrD[24:20]),
		.Funct3D(InstrD[14:12]),
		.IntDivE(IntDivE),
		.InstrD(InstrD),
		.StallE(StallE),
		.StallM(StallM),
		.StallW(StallW),
		.FlushE(FlushE),
		.FlushM(FlushM),
		.FlushW(FlushW),
		.FRM_REGW(FRM_REGW),
		.STATUS_FS(STATUS_FS),
		.FDivBusyE(FDivBusyE),
		.reset(reset),
		.clk(clk),
		.FRegWriteE(FRegWriteE),
		.FRegWriteM(FRegWriteM),
		.FRegWriteW(FRegWriteW),
		.ZfaE(ZfaE),
		.ZfaM(ZfaM),
		.ZfaFRoundNXE(ZfaFRoundNXE),
		.FrmE(FrmE),
		.FrmM(FrmM),
		.FmtE(FmtE),
		.FmtM(FmtM),
		.FDivStartE(FDivStartE),
		.IDivStartE(IDivStartE),
		.FWriteIntE(FWriteIntE),
		.FCvtIntE(FCvtIntE),
		.FWriteIntM(FWriteIntM),
		.OpCtrlE(OpCtrlE),
		.OpCtrlM(OpCtrlM),
		.FpLoadStoreM(FpLoadStoreM),
		.IllegalFPUInstrD(IllegalFPUInstrD),
		.XEnD(XEnD),
		.YEnD(YEnD),
		.ZEnD(ZEnD),
		.XEnE(XEnE),
		.YEnE(YEnE),
		.ZEnE(ZEnE),
		.FResSelE(FResSelE),
		.FResSelM(FResSelM),
		.FResSelW(FResSelW),
		.FPUActiveE(FPUActiveE),
		.PostProcSelE(PostProcSelE),
		.PostProcSelM(PostProcSelM),
		.FCvtIntW(FCvtIntW),
		.Adr1D(Adr1D),
		.Adr2D(Adr2D),
		.Adr3D(Adr3D),
		.Adr1E(Adr1E),
		.Adr2E(Adr2E),
		.Adr3E(Adr3E)
	);
	fregfile #(.FLEN($signed(P[901-:32]))) fregfile(
		.clk(clk),
		.reset(reset),
		.we4(FRegWriteW),
		.a1(InstrD[19:15]),
		.a2(InstrD[24:20]),
		.a3(InstrD[31:27]),
		.a4(RdW),
		.wd4(FResultW),
		.rd1(FRD1D),
		.rd2(FRD2D),
		.rd3(FRD3D)
	);
	flopenrc #(.WIDTH($signed(P[901-:32]))) DEReg1(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(FRD1D),
		.q(FRD1E)
	);
	flopenrc #(.WIDTH($signed(P[901-:32]))) DEReg2(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(FRD2D),
		.q(FRD2E)
	);
	flopenrc #(.WIDTH($signed(P[901-:32]))) DEReg3(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(FRD3D),
		.q(FRD3E)
	);
	fhazard fhazard(
		.Adr1D(Adr1D),
		.Adr2D(Adr2D),
		.Adr3D(Adr3D),
		.Adr1E(Adr1E),
		.Adr2E(Adr2E),
		.Adr3E(Adr3E),
		.FRegWriteE(FRegWriteE),
		.FRegWriteM(FRegWriteM),
		.FRegWriteW(FRegWriteW),
		.RdE(RdE),
		.RdM(RdM),
		.RdW(RdW),
		.FResSelM(FResSelM),
		.XEnD(XEnD),
		.YEnD(YEnD),
		.ZEnD(ZEnD),
		.FPUStallD(FPUStallD),
		.ForwardXE(ForwardXE),
		.ForwardYE(ForwardYE),
		.ForwardZE(ForwardZE)
	);
	mux3 #(.WIDTH($signed(P[901-:32]))) fxemux(
		.d0(FRD1E),
		.d1(FResultW),
		.d2(PreFpResM),
		.s(ForwardXE),
		.y(XE)
	);
	mux3 #(.WIDTH($signed(P[901-:32]))) fyemux(
		.d0(FRD2E),
		.d1(FResultW),
		.d2(PreFpResM),
		.s(ForwardYE),
		.y(PreYE)
	);
	mux3 #(.WIDTH($signed(P[901-:32]))) fzemux(
		.d0(FRD3E),
		.d1(FResultW),
		.d2(PreFpResM),
		.s(ForwardZE),
		.y(PreZE)
	);
	function automatic signed [$signed(P[1097-:32]) - 1:0] sv2v_cast_CACF9_signed;
		input reg signed [$signed(P[1097-:32]) - 1:0] inp;
		sv2v_cast_CACF9_signed = inp;
	endfunction
	function automatic signed [$signed(P[1227-:32]) - 1:0] sv2v_cast_4FCCE_signed;
		input reg signed [$signed(P[1227-:32]) - 1:0] inp;
		sv2v_cast_4FCCE_signed = inp;
	endfunction
	function automatic signed [$signed(P[967-:32]) - 1:0] sv2v_cast_17AC2_signed;
		input reg signed [$signed(P[967-:32]) - 1:0] inp;
		sv2v_cast_17AC2_signed = inp;
	endfunction
	function automatic signed [$signed(P[805-:32]) - 1:0] sv2v_cast_C2987_signed;
		input reg signed [$signed(P[805-:32]) - 1:0] inp;
		sv2v_cast_C2987_signed = inp;
	endfunction
	function automatic signed [$signed(P[611-:32]) - 1:0] sv2v_cast_C55D7_signed;
		input reg signed [$signed(P[611-:32]) - 1:0] inp;
		sv2v_cast_C55D7_signed = inp;
	endfunction
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk1
			assign BoxedOneE = {2'b00, {$signed(P[837-:32]) - 1 {1'b1}}, sv2v_cast_C2987_signed(0)};
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk1
			mux2 #(.WIDTH($signed(P[901-:32]))) fonemux(
				.d0({{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 2'b00, {$signed(P[643-:32]) - 1 {1'b1}}, sv2v_cast_C55D7_signed(0)}),
				.d1({2'b00, {$signed(P[837-:32]) - 1 {1'b1}}, sv2v_cast_C2987_signed(0)}),
				.s(FmtE),
				.y(BoxedOneE)
			);
		end
		else if (($signed(P[739-:32]) == 3) | ($signed(P[739-:32]) == 4)) begin : genblk1
			mux4 #(.WIDTH($signed(P[901-:32]))) fonemux(
				.d0({{$signed(P[901-:32]) - $signed(P[1161-:32]) {1'b1}}, 2'b00, {$signed(P[1129-:32]) - 1 {1'b1}}, sv2v_cast_CACF9_signed(0)}),
				.d1({{$signed(P[901-:32]) - $signed(P[1291-:32]) {1'b1}}, 2'b00, {$signed(P[1259-:32]) - 1 {1'b1}}, sv2v_cast_4FCCE_signed(0)}),
				.d2({{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, 2'b00, {$signed(P[999-:32]) - 1 {1'b1}}, sv2v_cast_17AC2_signed(0)}),
				.d3({2'b00, {$signed(P[837-:32]) - 1 {1'b1}}, sv2v_cast_C2987_signed(0)}),
				.s(FmtE),
				.y(BoxedOneE)
			);
		end
	endgenerate
	assign FmaAddSubE = (OpCtrlE[2] & OpCtrlE[1]) & (PostProcSelE == 2'b10);
	mux2 #(.WIDTH($signed(P[901-:32]))) fyaddmux(
		.d0(PreYE),
		.d1(BoxedOneE),
		.s(FmaAddSubE),
		.y(YE)
	);
	function automatic signed [$signed(P[901-:32]) - 1:0] sv2v_cast_7604C_signed;
		input reg signed [$signed(P[901-:32]) - 1:0] inp;
		sv2v_cast_7604C_signed = inp;
	endfunction
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk2
			assign BoxedZeroE = 1'sb0;
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk2
			mux2 #(.WIDTH($signed(P[901-:32]))) fmulzeromux(
				.d0({{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, {$signed(P[675-:32]) {1'b0}}}),
				.d1(sv2v_cast_7604C_signed(0)),
				.s(FmtE),
				.y(BoxedZeroE)
			);
		end
		else if (($signed(P[739-:32]) == 3) | ($signed(P[739-:32]) == 4)) begin : genblk2
			mux4 #(.WIDTH($signed(P[901-:32]))) fmulzeromux(
				.d0({{$signed(P[901-:32]) - $signed(P[1161-:32]) {1'b1}}, {$signed(P[1161-:32]) {1'b0}}}),
				.d1({{$signed(P[901-:32]) - $signed(P[1291-:32]) {1'b1}}, {$signed(P[1291-:32]) {1'b0}}}),
				.d2({{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, {$signed(P[1031-:32]) {1'b0}}}),
				.d3(sv2v_cast_7604C_signed(0)),
				.s(FmtE),
				.y(BoxedZeroE)
			);
		end
	endgenerate
	assign FmaZSelE = {OpCtrlE[2] & OpCtrlE[1], OpCtrlE[2] & ~OpCtrlE[1]};
	mux3 #(.WIDTH($signed(P[901-:32]))) fzmulmux(
		.d0(PreZE),
		.d1(BoxedZeroE),
		.d2(PreYE),
		.s(FmaZSelE),
		.y(ZE)
	);
	unpack #(.P(P)) unpack(
		.X(XE),
		.Y(YE),
		.Z(ZE),
		.Fmt(FmtE),
		.Xs(XsE),
		.Ys(YsE),
		.Zs(ZsE),
		.Xe(XeE),
		.Ye(YeE),
		.Ze(ZeE),
		.Xm(XmE),
		.Ym(YmE),
		.Zm(ZmE),
		.YEn(YEnE),
		.FPUActive(FPUActiveE),
		.XNaN(XNaNE),
		.YNaN(YNaNE),
		.ZNaN(ZNaNE),
		.XSNaN(XSNaNE),
		.XEn(XEnE),
		.YSNaN(YSNaNE),
		.ZSNaN(ZSNaNE),
		.XSubnorm(XSubnormE),
		.XZero(XZeroE),
		.YZero(YZeroE),
		.ZZero(ZZeroE),
		.XInf(XInfE),
		.YInf(YInfE),
		.ZEn(ZEnE),
		.ZInf(ZInfE),
		.XExpMax(XExpMaxE),
		.XPostBox(XPostBoxE),
		.Bias(BiasE),
		.Nf(NfE)
	);
	fma #(.P(P)) fma(
		.Xs(XsE),
		.Ys(YsE),
		.Zs(ZsE),
		.Xe(XeE),
		.Ye(YeE),
		.Ze(ZeE),
		.Xm(XmE),
		.Ym(YmE),
		.Zm(ZmE),
		.XZero(XZeroE),
		.YZero(YZeroE),
		.ZZero(ZZeroE),
		.OpCtrl(OpCtrlE),
		.As(AsE),
		.Ps(PsE),
		.Ss(SsE),
		.Se(SeE),
		.Sm(SmE),
		.InvA(InvAE),
		.SCnt(SCntE),
		.ASticky(FmaAStickyE)
	);
	fdivsqrt #(.P(P)) fdivsqrt(
		.clk(clk),
		.reset(reset),
		.FmtE(FmtE),
		.XmE(XmE),
		.YmE(YmE),
		.XeE(XeE),
		.YeE(YeE),
		.SqrtE(OpCtrlE[0]),
		.SqrtM(OpCtrlM[0]),
		.XInfE(XInfE),
		.YInfE(YInfE),
		.XZeroE(XZeroE),
		.YZeroE(YZeroE),
		.XNaNE(XNaNE),
		.YNaNE(YNaNE),
		.BiasE(BiasE),
		.NfE(NfE),
		.FDivStartE(FDivStartE),
		.IDivStartE(IDivStartE),
		.XsE(XsE),
		.ForwardedSrcAE(ForwardedSrcAE),
		.ForwardedSrcBE(ForwardedSrcBE),
		.Funct3E(Funct3E),
		.Funct3M(Funct3M),
		.IntDivE(IntDivE),
		.W64E(W64E),
		.StallM(StallM),
		.FlushE(FlushE),
		.DivStickyM(DivStickyM),
		.FDivBusyE(FDivBusyE),
		.IFDivStartE(IFDivStartE),
		.FDivDoneE(FDivDoneE),
		.UeM(UeM),
		.UmM(UmM),
		.FIntDivResultM(FIntDivResultM)
	);
	fcmp #(.P(P)) fcmp(
		.Fmt(FmtE),
		.OpCtrl(OpCtrlE),
		.Zfa(ZfaE),
		.Xs(XsE),
		.Ys(YsE),
		.Xe(XeE),
		.Ye(YeE),
		.Xm(XmE),
		.Ym(YmE),
		.XZero(XZeroE),
		.YZero(YZeroE),
		.XNaN(XNaNE),
		.YNaN(YNaNE),
		.XSNaN(XSNaNE),
		.YSNaN(YSNaNE),
		.X(XE),
		.Y(YE),
		.CmpNV(CmpNVE),
		.CmpFpRes(CmpFpResE),
		.CmpIntRes(CmpIntResE)
	);
	fsgninj #(.P(P)) fsgninj(
		.OpCtrl(OpCtrlE[1:0]),
		.Xs(XsE),
		.Ys(YsE),
		.X(XPostBoxE),
		.Fmt(FmtE),
		.SgnRes(SgnResE)
	);
	fclassify #(.P(P)) fclassify(
		.Xs(XsE),
		.XSubnorm(XSubnormE),
		.XZero(XZeroE),
		.XNaN(XNaNE),
		.XInf(XInfE),
		.XSNaN(XSNaNE),
		.ClassRes(ClassResE)
	);
	fcvt #(.P(P)) fcvt(
		.Xs(XsE),
		.Xe(XeE),
		.Xm(XmE),
		.Int(ForwardedSrcAE),
		.OpCtrl(OpCtrlE),
		.ToInt(FWriteIntE),
		.XZero(XZeroE),
		.Fmt(FmtE),
		.Ce(CeE),
		.ShiftAmt(CvtShiftAmtE),
		.ResSubnormUf(CvtResSubnormUfE),
		.Cs(CsE),
		.IntZero(IntZeroE),
		.LzcIn(CvtLzcInE)
	);
	generate
		if (P[4069]) begin : Zfa
			wire [4:0] Rs1E;
			wire [1:0] Fmt2E;
			wire [$signed(P[901-:32]) - 1:0] FRoundE;
			wire [$signed(P[901-:32]) - 1:0] FliResE;
			fround #(.P(P)) fround(
				.Xs(XsE),
				.Xe(XeE),
				.Xm(XmE),
				.XNaN(XNaNE),
				.XSNaN(XSNaNE),
				.Fmt(FmtE),
				.Frm(FrmE),
				.Nf(NfE),
				.ZfaFRoundNX(ZfaFRoundNXE),
				.FRound(FRoundE),
				.FRoundNV(FRoundNVE),
				.FRoundNX(FRoundNXE)
			);
			flopenrc #(.WIDTH(5)) Rs1EReg(
				.clk(clk),
				.reset(reset),
				.clear(FlushE),
				.en(~StallE),
				.d(InstrD[19:15]),
				.q(Rs1E)
			);
			flopenrc #(.WIDTH(2)) Fmt2EReg(
				.clk(clk),
				.reset(reset),
				.clear(FlushE),
				.en(~StallE),
				.d(InstrD[26:25]),
				.q(Fmt2E)
			);
			fli #(.P(P)) fli(
				.Rs1(Rs1E),
				.Fmt(Fmt2E),
				.Imm(FliResE)
			);
			mux2 #(.WIDTH($signed(P[901-:32]))) ZfaResMux(
				.d0(FRoundE),
				.d1(FliResE),
				.s(OpCtrlE[0]),
				.y(ZfaResE)
			);
		end
		else begin : genblk3
			assign {FRoundNXE, FRoundNVE} = 1'sb0;
			assign ZfaResE = 1'sbx;
		end
		if ($signed(P[739-:32]) == 1) begin : genblk4
			if ($signed(P[901-:32]) >= $signed(P[4216-:32])) begin : genblk1
				assign PreIntSrcE = {{$signed(P[901-:32]) - $signed(P[4216-:32]) {1'b1}}, ForwardedSrcAE};
			end
			else begin : genblk1
				assign PreIntSrcE = ForwardedSrcAE[$signed(P[901-:32]) - 1:0];
			end
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk4
			if ($signed(P[901-:32]) >= $signed(P[4216-:32])) begin : genblk1
				mux2 #(.WIDTH($signed(P[901-:32]))) SrcAMux(
					.d0({{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, ForwardedSrcAE[$signed(P[675-:32]) - 1:0]}),
					.d1({{$signed(P[901-:32]) - $signed(P[4216-:32]) {1'b1}}, ForwardedSrcAE}),
					.s(FmtE),
					.y(PreIntSrcE)
				);
			end
			else begin : genblk1
				mux2 #(.WIDTH($signed(P[901-:32]))) SrcAMux(
					.d0({{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, ForwardedSrcAE[$signed(P[675-:32]) - 1:0]}),
					.d1(ForwardedSrcAE[$signed(P[901-:32]) - 1:0]),
					.s(FmtE),
					.y(PreIntSrcE)
				);
			end
		end
		else if (($signed(P[739-:32]) == 3) | ($signed(P[739-:32]) == 4)) begin : genblk4
			localparam XD_LEN = ($signed(P[1291-:32]) < $signed(P[4216-:32]) ? $signed(P[1291-:32]) : $signed(P[4216-:32]));
			mux3 #(.WIDTH($signed(P[901-:32]))) SrcAMux(
				.d0({{$signed(P[901-:32]) - $signed(P[1161-:32]) {1'b1}}, ForwardedSrcAE[$signed(P[1161-:32]) - 1:0]}),
				.d1({{$signed(P[901-:32]) - XD_LEN {1'b1}}, ForwardedSrcAE[XD_LEN - 1:0]}),
				.d2({{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, ForwardedSrcAE[$signed(P[1031-:32]) - 1:0]}),
				.s(FmtE),
				.y(PreIntSrcE)
			);
		end
		if (P[4069] & ($signed(P[901-:32]) == (2 * $signed(P[4216-:32])))) begin : genblk5
			assign IntSrcE = (ZfaE ? {ForwardedSrcBE, ForwardedSrcAE} : PreIntSrcE);
		end
		else begin : genblk5
			assign IntSrcE = PreIntSrcE;
		end
	endgenerate
	mux4 #(.WIDTH($signed(P[901-:32]))) FResMux(
		.d0(SgnResE),
		.d1(IntSrcE),
		.d2(CmpFpResE),
		.d3(ZfaResE),
		.s({OpCtrlE[2], &OpCtrlE[1:0] | ((OpCtrlE == 3'b100) & ZfaE)}),
		.y(PreFpResE)
	);
	assign PreNVE = (CmpNVE & (OpCtrlE[2] | FWriteIntE)) | ((FRoundNVE & (OpCtrlE == 3'b100)) & ZfaE);
	assign PreNXE = FRoundNXE & (OpCtrlE == 3'b100);
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk6
			assign mvsgn = XE[$signed(P[901-:32]) - 1];
			assign SgnExtXE = XE;
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk6
			mux2 #(.WIDTH(1)) sgnmux(
				.d0(XE[$signed(P[675-:32]) - 1]),
				.d1(XE[$signed(P[901-:32]) - 1]),
				.s(FmtE),
				.y(mvsgn)
			);
			mux2 #(.WIDTH($signed(P[901-:32]))) sgnextmux(
				.d0({{$signed(P[901-:32]) - $signed(P[675-:32]) {mvsgn}}, XE[$signed(P[675-:32]) - 1:0]}),
				.d1(XE),
				.s(FmtE),
				.y(SgnExtXE)
			);
		end
		else if (($signed(P[739-:32]) == 3) | ($signed(P[739-:32]) == 4)) begin : genblk6
			mux4 #(.WIDTH(1)) sgnmux(
				.d0(XE[$signed(P[1161-:32]) - 1]),
				.d1(XE[$signed(P[1291-:32]) - 1]),
				.d2(XE[$signed(P[1031-:32]) - 1]),
				.d3(XE[$signed(P[383-:32]) - 1]),
				.s(FmtE),
				.y(mvsgn)
			);
			mux3 #(.WIDTH($signed(P[901-:32]))) sgnextmux(
				.d0({{$signed(P[901-:32]) - $signed(P[1161-:32]) {mvsgn}}, XE[$signed(P[1161-:32]) - 1:0]}),
				.d1({{$signed(P[901-:32]) - $signed(P[1291-:32]) {mvsgn}}, XE[$signed(P[1291-:32]) - 1:0]}),
				.d2({{$signed(P[901-:32]) - $signed(P[1031-:32]) {mvsgn}}, XE[$signed(P[1031-:32]) - 1:0]}),
				.s(FmtE),
				.y(SgnExtXE)
			);
		end
		if ($signed(P[901-:32]) >= (2 * $signed(P[4216-:32]))) begin : genblk7
			if (P[4069]) begin : genblk1
				assign IntSrcXE = (ZfaE ? XE[(2 * $signed(P[4216-:32])) - 1:$signed(P[4216-:32])] : SgnExtXE[$signed(P[4216-:32]) - 1:0]);
			end
			else begin : genblk1
				assign IntSrcXE = SgnExtXE[$signed(P[4216-:32]) - 1:0];
			end
		end
		else begin : genblk7
			assign IntSrcXE = {{$signed(P[4216-:32]) - $signed(P[901-:32]) {mvsgn}}, SgnExtXE};
		end
	endgenerate
	mux3 #(.WIDTH($signed(P[4216-:32]))) IntResMux(
		.d0(ClassResE),
		.d1(IntSrcXE),
		.d2(CmpIntResE),
		.s({~FResSelE[1], FResSelE[0]}),
		.y(FIntResE)
	);
	assign StallUnpackedM = StallM | ((FDivBusyE & ~IFDivStartE) | FDivDoneE);
	flopenrc #(.WIDTH($signed(P[805-:32]) + 1)) EMFpReg2(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(XmE),
		.q(XmM)
	);
	flopenrc #(.WIDTH($signed(P[805-:32]) + 1)) EMFpReg3(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(YmE),
		.q(YmM)
	);
	flopenrc #(.WIDTH($signed(P[901-:32]))) EMFpReg4(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d({ZeE, ZmE}),
		.q({ZeM, ZmM})
	);
	flopenrc #(.WIDTH($signed(P[4216-:32]))) EMFpReg6(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(FIntResE),
		.q(FIntResM)
	);
	flopenrc #(.WIDTH($signed(P[901-:32]))) EMFpReg7(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(PreFpResE),
		.q(PreFpResM)
	);
	flopenr #(.WIDTH(13)) EMFpReg5(
		.clk(clk),
		.reset(reset),
		.en(~StallUnpackedM),
		.d({XsE, YsE, XZeroE, YZeroE, XInfE, YInfE, ZInfE, XNaNE, YNaNE, ZNaNE, XSNaNE, YSNaNE, ZSNaNE}),
		.q({XsM, YsM, XZeroM, YZeroM, XInfM, YInfM, ZInfM, XNaNM, YNaNM, ZNaNM, XSNaNM, YSNaNM, ZSNaNM})
	);
	flopenrc #(.WIDTH(2)) EMRegCmpFlg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d({PreNVE, PreNXE}),
		.q({PreNVM, PreNXM})
	);
	flopenrc #(.WIDTH($signed(P[255-:32]))) EMRegFma2(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(SmE),
		.q(SmM)
	);
	flopenrc #(.WIDTH(($clog2($signed(P[255-:32]) + 1) + 7) + $signed(P[837-:32]))) EMRegFma4(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d({FmaAStickyE, InvAE, SCntE, AsE, PsE, SsE, SeE}),
		.q({FmaAStickyM, InvAM, SCntM, AsM, PsM, SsM, SeM})
	);
	flopenrc #(.WIDTH((($signed(P[837-:32]) + $signed(P[351-:32])) + $signed(P[415-:32])) + 4)) EMRegCvt(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d({CeE, CvtShiftAmtE, CvtResSubnormUfE, CsE, IntZeroE, CvtLzcInE}),
		.q({CeM, CvtShiftAmtM, CvtResSubnormUfM, CsM, IntZeroM, CvtLzcInM})
	);
	flopenrc #(.WIDTH($signed(P[901-:32]))) FWriteDataMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(YE),
		.q(FWriteDataM)
	);
	postprocess #(.P(P)) postprocess(
		.Xs(XsM),
		.Ys(YsM),
		.Xm(XmM),
		.Ym(YmM),
		.Zm(ZmM),
		.Frm(FrmM),
		.Fmt(FmtM),
		.FmaASticky(FmaAStickyM),
		.XZero(XZeroM),
		.YZero(YZeroM),
		.XInf(XInfM),
		.YInf(YInfM),
		.DivUm(UmM),
		.FmaSs(SsM),
		.ZInf(ZInfM),
		.XNaN(XNaNM),
		.YNaN(YNaNM),
		.ZNaN(ZNaNM),
		.XSNaN(XSNaNM),
		.YSNaN(YSNaNM),
		.ZSNaN(ZSNaNM),
		.FmaSm(SmM),
		.DivUe(UeM),
		.FmaAs(AsM),
		.FmaPs(PsM),
		.OpCtrl(OpCtrlM),
		.FmaSCnt(SCntM),
		.FmaSe(SeM),
		.CvtCe(CeM),
		.CvtResSubnormUf(CvtResSubnormUfM),
		.CvtShiftAmt(CvtShiftAmtM),
		.CvtCs(CsM),
		.ToInt(FWriteIntM),
		.Zfa(ZfaM),
		.DivSticky(DivStickyM),
		.CvtLzcIn(CvtLzcInM),
		.IntZero(IntZeroM),
		.PostProcSel(PostProcSelM),
		.PostProcRes(PostProcResM),
		.PostProcFlg(PostProcFlgM),
		.FCvtIntRes(FCvtIntResM)
	);
	mux2 #(.WIDTH(5)) FPUFlgMux(
		.d0({PreNVM, 3'b000, PreNXM}),
		.d1(PostProcFlgM),
		.s(FResSelM == 2'b01),
		.y(SetFflagsM)
	);
	mux2 #(.WIDTH($signed(P[901-:32]))) FPUResMux(
		.d0(PreFpResM),
		.d1(PostProcResM),
		.s(FResSelM[0]),
		.y(FpResM)
	);
	flopenrc #(.WIDTH($signed(P[901-:32]))) MWRegFp(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(FpResM),
		.q(FpResW)
	);
	flopenrc #(.WIDTH($signed(P[4216-:32]))) MWRegIntCvtRes(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(FCvtIntResM),
		.q(FCvtIntResW)
	);
	flopenrc #(.WIDTH($signed(P[4216-:32]))) MWRegIntDivRes(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(FIntDivResultM),
		.q(FIntDivResultW)
	);
	mux2 #(.WIDTH($signed(P[901-:32]))) FResultMux(
		.d0(FpResW),
		.d1(ReadDataW),
		.s(FResSelW[1]),
		.y(FResultW)
	);
endmodule
module fregfile (
	clk,
	reset,
	we4,
	a1,
	a2,
	a3,
	a4,
	wd4,
	rd1,
	rd2,
	rd3
);
	parameter FLEN = 0;
	input wire clk;
	input wire reset;
	input wire we4;
	input wire [4:0] a1;
	input wire [4:0] a2;
	input wire [4:0] a3;
	input wire [4:0] a4;
	input wire [FLEN - 1:0] wd4;
	output wire [FLEN - 1:0] rd1;
	output wire [FLEN - 1:0] rd2;
	output wire [FLEN - 1:0] rd3;
	reg [FLEN - 1:0] rf [31:0];
	integer i;
	always @(negedge clk)
		if (reset)
			for (i = 0; i < 32; i = i + 1)
				rf[i] <= 1'sb0;
		else if (we4)
			rf[a4] <= wd4;
	assign rd1 = rf[a1];
	assign rd2 = rf[a2];
	assign rd3 = rf[a3];
endmodule
module fround (
	Xs,
	Xe,
	Xm,
	XNaN,
	XSNaN,
	Fmt,
	Frm,
	Nf,
	ZfaFRoundNX,
	FRound,
	FRoundNV,
	FRoundNX
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire Xs;
	input wire [$signed(P[837-:32]) - 1:0] Xe;
	input wire [$signed(P[805-:32]):0] Xm;
	input wire XNaN;
	input wire XSNaN;
	input wire [$signed(P[707-:32]) - 1:0] Fmt;
	input wire [2:0] Frm;
	input wire [$signed(P[869-:32]) - 1:0] Nf;
	input wire ZfaFRoundNX;
	output wire [$signed(P[901-:32]) - 1:0] FRound;
	output wire FRoundNV;
	output wire FRoundNX;
	wire [$signed(P[837-:32]) - 1:0] E;
	wire [$signed(P[837-:32]) - 1:0] Xep1;
	wire [$signed(P[805-:32]):0] IMask;
	wire [$signed(P[805-:32]):0] Tmasknonneg;
	wire [$signed(P[805-:32]):0] Tmaskneg;
	wire [$signed(P[805-:32]):0] Tmask;
	wire [$signed(P[805-:32]):0] HotE;
	wire [$signed(P[805-:32]):0] HotEP1;
	wire [$signed(P[805-:32]):0] Trunc;
	wire [$signed(P[805-:32]):0] Rnd;
	reg [$signed(P[901-:32]) - 1:0] W;
	wire Elt0;
	wire Eeqm1;
	wire Lnonneg;
	wire Lp;
	wire Rnonneg;
	wire Rp;
	wire Tp;
	reg RoundUp;
	wire Two;
	wire EgeNf;
	assign E = Xe - P[739 + $signed(P[837-:32]):740];
	assign Xep1 = Xe + 1'b1;
	assign Elt0 = E[$signed(P[837-:32]) - 1];
	assign Eeqm1 = $signed(E) == -1;
	assign IMask = $signed({1'b1, {$signed(P[805-:32]) {1'b0}}}) >>> E;
	assign Tmasknonneg = ~IMask >>> 1'b1;
	assign HotE = IMask & ~(IMask << 1'b1);
	assign HotEP1 = HotE >> 1'b1;
	assign Lnonneg = |(Xm & HotE);
	assign Rnonneg = |(Xm & HotEP1);
	assign Trunc = Xm & IMask;
	assign {Two, Rnd} = Trunc + HotE;
	mux2 #(.WIDTH(1)) Lmux(
		.d0(Lnonneg),
		.d1(1'b0),
		.s(Elt0),
		.y(Lp)
	);
	mux2 #(.WIDTH(1)) Rmux(
		.d0(Rnonneg),
		.d1(Eeqm1),
		.s(Elt0),
		.y(Rp)
	);
	assign Tmaskneg = {~Eeqm1, {$signed(P[805-:32]) {1'b1}}};
	mux2 #(.WIDTH($signed(P[805-:32]) + 1)) Tmaskmux(
		.d0(Tmasknonneg),
		.d1(Tmaskneg),
		.s(Elt0),
		.y(Tmask)
	);
	assign Tp = |(Xm & Tmask);
	assign EgeNf = (E >= Nf) & Xe[$signed(P[837-:32]) - 1];
	always @(*) begin
		if (_sv2v_0)
			;
		case (Frm)
			3'b000: RoundUp = Rp & (Lp | Tp);
			3'b001: RoundUp = 0;
			3'b010: RoundUp = Xs & (Rp | Tp);
			3'b011: RoundUp = ~Xs & (Rp | Tp);
			3'b100: RoundUp = Rp;
			default: RoundUp = 0;
		endcase
		if (XNaN)
			W = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, {$signed(P[805-:32]) - 1 {1'b0}}};
		else if (EgeNf)
			W = {Xs, Xe, Xm[$signed(P[805-:32]) - 1:0]};
		else if (Elt0) begin
			if (RoundUp)
				W = {Xs, P[739 + $signed(P[837-:32]):740], {$signed(P[805-:32]) {1'b0}}};
			else
				W = {Xs, {$signed(P[901-:32]) - 1 {1'b0}}};
		end
		else if (RoundUp & Two)
			W = {Xs, Xep1, {$signed(P[805-:32]) {1'b0}}};
		else if (RoundUp)
			W = {Xs, Xe, Rnd[$signed(P[805-:32]) - 1:0]};
		else
			W = {Xs, Xe, Trunc[$signed(P[805-:32]) - 1:0]};
	end
	packoutput #(.P(P)) packoutput(
		.Unpacked(W),
		.Fmt(Fmt),
		.Packed(FRound)
	);
	assign FRoundNV = XSNaN;
	assign FRoundNX = ((ZfaFRoundNX & ~EgeNf) & (Rp | Tp)) & ~XNaN;
	initial _sv2v_0 = 0;
endmodule
module fsgninj (
	Xs,
	Ys,
	X,
	Fmt,
	OpCtrl,
	SgnRes
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire Xs;
	input wire Ys;
	input wire [$signed(P[901-:32]) - 1:0] X;
	input wire [$signed(P[707-:32]) - 1:0] Fmt;
	input wire [1:0] OpCtrl;
	output wire [$signed(P[901-:32]) - 1:0] SgnRes;
	wire ResSgn;
	assign ResSgn = (OpCtrl[1] ? Xs : OpCtrl[0]) ^ Ys;
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk1
			assign SgnRes = {ResSgn, X[$signed(P[901-:32]) - 2:0]};
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk1
			assign SgnRes = {~Fmt | ResSgn, X[$signed(P[901-:32]) - 2:$signed(P[675-:32])], (Fmt ? X[$signed(P[675-:32]) - 1] : ResSgn), X[$signed(P[675-:32]) - 2:0]};
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk1
			reg [2:0] SgnBits;
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					P[773-:2]: SgnBits = {ResSgn, X[$signed(P[675-:32]) - 1], X[$signed(P[545-:32]) - 1]};
					P[579-:2]: SgnBits = {1'b1, ResSgn, X[$signed(P[545-:32]) - 1]};
					P[449-:2]: SgnBits = {2'b11, ResSgn};
					default: SgnBits = {3 {1'bx}};
				endcase
			end
			assign SgnRes = {SgnBits[2], X[$signed(P[901-:32]) - 2:$signed(P[675-:32])], SgnBits[1], X[$signed(P[675-:32]) - 2:$signed(P[545-:32])], SgnBits[0], X[$signed(P[545-:32]) - 2:0]};
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk1
			reg [3:0] SgnBits;
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					P[1293-:2]: SgnBits = {ResSgn, X[$signed(P[1291-:32]) - 1], X[$signed(P[1161-:32]) - 1], X[$signed(P[1031-:32]) - 1]};
					P[1163-:2]: SgnBits = {1'b1, ResSgn, X[$signed(P[1161-:32]) - 1], X[$signed(P[1031-:32]) - 1]};
					P[1033-:2]: SgnBits = {2'b11, ResSgn, X[$signed(P[1031-:32]) - 1]};
					P[903-:2]: SgnBits = {3'b111, ResSgn};
				endcase
			end
			assign SgnRes = {SgnBits[3], X[$signed(P[1421-:32]) - 2:$signed(P[1291-:32])], SgnBits[2], X[$signed(P[1291-:32]) - 2:$signed(P[1161-:32])], SgnBits[1], X[$signed(P[1161-:32]) - 2:$signed(P[1031-:32])], SgnBits[0], X[$signed(P[1031-:32]) - 2:0]};
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module packoutput (
	Unpacked,
	Fmt,
	Packed
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[901-:32]) - 1:0] Unpacked;
	input wire [$signed(P[707-:32]) - 1:0] Fmt;
	output reg [$signed(P[901-:32]) - 1:0] Packed;
	wire Sign;
	reg [$signed(P[643-:32]) - 1:0] Exp1;
	reg [$signed(P[611-:32]) - 1:0] Fract1;
	reg [$signed(P[513-:32]) - 1:0] Exp2;
	reg [$signed(P[481-:32]) - 1:0] Fract2;
	reg [$signed(P[999-:32]) - 1:0] Exp3;
	reg [$signed(P[967-:32]) - 1:0] Fract3;
	assign Sign = Unpacked[$signed(P[901-:32]) - 1];
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk1
			wire [$signed(P[901-:32]):1] sv2v_tmp_98EA2;
			assign sv2v_tmp_98EA2 = Unpacked;
			always @(*) Packed = sv2v_tmp_98EA2;
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				{Exp1, Fract1} = 1'sb0;
				case (Fmt)
					1'b1: Packed = Unpacked;
					1'b0: begin
						Exp1 = {Unpacked[$signed(P[901-:32]) - 2], Unpacked[($signed(P[805-:32]) + $signed(P[643-:32])) - 2:$signed(P[805-:32])]};
						Fract1 = Unpacked[$signed(P[805-:32]) - 1:$signed(P[805-:32]) - $signed(P[611-:32])];
						Packed = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, Sign, Exp1, Fract1};
					end
				endcase
			end
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				{Exp1, Fract1, Exp2, Fract2} = 1'sb0;
				case (Fmt)
					P[773-:2]: Packed = Unpacked;
					P[579-:2]: begin
						Exp1 = {Unpacked[$signed(P[901-:32]) - 2], Unpacked[($signed(P[805-:32]) + $signed(P[643-:32])) - 2:$signed(P[805-:32])]};
						Fract1 = Unpacked[$signed(P[805-:32]) - 1:$signed(P[805-:32]) - $signed(P[611-:32])];
						Packed = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, Sign, Exp1, Fract1};
					end
					P[449-:2]: begin
						Exp2 = {Unpacked[$signed(P[901-:32]) - 2], Unpacked[($signed(P[805-:32]) + $signed(P[513-:32])) - 2:$signed(P[805-:32])]};
						Fract2 = Unpacked[$signed(P[805-:32]) - 1:$signed(P[805-:32]) - $signed(P[481-:32])];
						Packed = {{$signed(P[901-:32]) - $signed(P[545-:32]) {1'b1}}, Sign, Exp2, Fract2};
					end
					default: Packed = 1'sbx;
				endcase
			end
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				{Exp1, Fract1, Exp2, Fract2, Exp3, Fract3} = 1'sb0;
				case (Fmt)
					2'h3: Packed = Unpacked;
					2'h1: begin
						Exp1 = {Unpacked[$signed(P[901-:32]) - 2], Unpacked[($signed(P[805-:32]) + $signed(P[643-:32])) - 2:$signed(P[805-:32])]};
						Fract1 = Unpacked[$signed(P[805-:32]) - 1:$signed(P[805-:32]) - $signed(P[611-:32])];
						Packed = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, Sign, Exp1, Fract1};
					end
					2'h0: begin
						Exp2 = {Unpacked[$signed(P[901-:32]) - 2], Unpacked[($signed(P[805-:32]) + $signed(P[513-:32])) - 2:$signed(P[805-:32])]};
						Fract2 = Unpacked[$signed(P[805-:32]) - 1:$signed(P[805-:32]) - $signed(P[481-:32])];
						Packed = {{$signed(P[901-:32]) - $signed(P[545-:32]) {1'b1}}, Sign, Exp2, Fract2};
					end
					2'h2: begin
						Exp3 = {Unpacked[$signed(P[901-:32]) - 2], Unpacked[($signed(P[805-:32]) + $signed(P[999-:32])) - 2:$signed(P[805-:32])]};
						Fract3 = Unpacked[$signed(P[805-:32]) - 1:$signed(P[805-:32]) - $signed(P[967-:32])];
						Packed = {{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, Sign, Exp3, Fract3};
					end
				endcase
			end
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module unpack (
	X,
	Y,
	Z,
	Fmt,
	XEn,
	YEn,
	ZEn,
	FPUActive,
	Xs,
	Ys,
	Zs,
	Xe,
	Ye,
	Ze,
	Xm,
	Ym,
	Zm,
	XNaN,
	YNaN,
	ZNaN,
	XSNaN,
	YSNaN,
	ZSNaN,
	XSubnorm,
	XZero,
	YZero,
	ZZero,
	XInf,
	YInf,
	ZInf,
	XExpMax,
	XPostBox,
	Bias,
	Nf
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[901-:32]) - 1:0] X;
	input wire [$signed(P[901-:32]) - 1:0] Y;
	input wire [$signed(P[901-:32]) - 1:0] Z;
	input wire [$signed(P[707-:32]) - 1:0] Fmt;
	input wire XEn;
	input wire YEn;
	input wire ZEn;
	input wire FPUActive;
	output wire Xs;
	output wire Ys;
	output wire Zs;
	output wire [$signed(P[837-:32]) - 1:0] Xe;
	output wire [$signed(P[837-:32]) - 1:0] Ye;
	output wire [$signed(P[837-:32]) - 1:0] Ze;
	output wire [$signed(P[805-:32]):0] Xm;
	output wire [$signed(P[805-:32]):0] Ym;
	output wire [$signed(P[805-:32]):0] Zm;
	output wire XNaN;
	output wire YNaN;
	output wire ZNaN;
	output wire XSNaN;
	output wire YSNaN;
	output wire ZSNaN;
	output wire XSubnorm;
	output wire XZero;
	output wire YZero;
	output wire ZZero;
	output wire XInf;
	output wire YInf;
	output wire ZInf;
	output wire XExpMax;
	output wire [$signed(P[901-:32]) - 1:0] XPostBox;
	output wire [$signed(P[837-:32]) - 2:0] Bias;
	output wire [$signed(P[869-:32]) - 1:0] Nf;
	wire YExpMax;
	wire ZExpMax;
	unpackinput #(.P(P)) unpackinputX(
		.A(X),
		.Fmt(Fmt),
		.Sgn(Xs),
		.Exp(Xe),
		.Man(Xm),
		.En(XEn),
		.FPUActive(FPUActive),
		.NaN(XNaN),
		.SNaN(XSNaN),
		.Zero(XZero),
		.Inf(XInf),
		.ExpMax(XExpMax),
		.Subnorm(XSubnorm),
		.PostBox(XPostBox)
	);
	unpackinput #(.P(P)) unpackinputY(
		.A(Y),
		.Fmt(Fmt),
		.Sgn(Ys),
		.Exp(Ye),
		.Man(Ym),
		.En(YEn),
		.FPUActive(FPUActive),
		.NaN(YNaN),
		.SNaN(YSNaN),
		.Zero(YZero),
		.Inf(YInf),
		.ExpMax(YExpMax),
		.Subnorm(),
		.PostBox()
	);
	unpackinput #(.P(P)) unpackinputZ(
		.A(Z),
		.Fmt(Fmt),
		.Sgn(Zs),
		.Exp(Ze),
		.Man(Zm),
		.En(ZEn),
		.FPUActive(FPUActive),
		.NaN(ZNaN),
		.SNaN(ZSNaN),
		.Zero(ZZero),
		.Inf(ZInf),
		.ExpMax(ZExpMax),
		.Subnorm(),
		.PostBox()
	);
	fmtparams #(.P(P)) fmtparams(
		.Fmt(Fmt),
		.Bias(Bias),
		.Nf(Nf)
	);
endmodule
module unpackinput (
	A,
	En,
	Fmt,
	FPUActive,
	Sgn,
	Exp,
	Man,
	NaN,
	SNaN,
	Zero,
	Inf,
	ExpMax,
	Subnorm,
	PostBox
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[901-:32]) - 1:0] A;
	input wire En;
	input wire [$signed(P[707-:32]) - 1:0] Fmt;
	input wire FPUActive;
	output reg Sgn;
	output reg [$signed(P[837-:32]) - 1:0] Exp;
	output wire [$signed(P[805-:32]):0] Man;
	output wire NaN;
	output wire SNaN;
	output wire Zero;
	output wire Inf;
	output reg ExpMax;
	output wire Subnorm;
	output reg [$signed(P[901-:32]) - 1:0] PostBox;
	reg [$signed(P[805-:32]) - 1:0] Frac;
	reg BadNaNBox;
	wire FracZero;
	reg ExpNonZero;
	wire [$signed(P[901-:32]) - 1:0] In;
	assign In = A & {$signed(P[901-:32]) {FPUActive}};
	function automatic signed [($signed(P[1357-:32]) - $signed(P[1227-:32])) - 1:0] sv2v_cast_FEE12_signed;
		input reg signed [($signed(P[1357-:32]) - $signed(P[1227-:32])) - 1:0] inp;
		sv2v_cast_FEE12_signed = inp;
	endfunction
	function automatic signed [($signed(P[1357-:32]) - $signed(P[1097-:32])) - 1:0] sv2v_cast_E94E5_signed;
		input reg signed [($signed(P[1357-:32]) - $signed(P[1097-:32])) - 1:0] inp;
		sv2v_cast_E94E5_signed = inp;
	endfunction
	function automatic signed [($signed(P[1357-:32]) - $signed(P[967-:32])) - 1:0] sv2v_cast_A7C1E_signed;
		input reg signed [($signed(P[1357-:32]) - $signed(P[967-:32])) - 1:0] inp;
		sv2v_cast_A7C1E_signed = inp;
	endfunction
	function automatic signed [($signed(P[805-:32]) - $signed(P[611-:32])) - 1:0] sv2v_cast_302A5_signed;
		input reg signed [($signed(P[805-:32]) - $signed(P[611-:32])) - 1:0] inp;
		sv2v_cast_302A5_signed = inp;
	endfunction
	function automatic signed [($signed(P[805-:32]) - $signed(P[481-:32])) - 1:0] sv2v_cast_8BF36_signed;
		input reg signed [($signed(P[805-:32]) - $signed(P[481-:32])) - 1:0] inp;
		sv2v_cast_8BF36_signed = inp;
	endfunction
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk1
			wire [1:1] sv2v_tmp_45FEF;
			assign sv2v_tmp_45FEF = 1'b0;
			always @(*) BadNaNBox = sv2v_tmp_45FEF;
			wire [1:1] sv2v_tmp_CA8B4;
			assign sv2v_tmp_CA8B4 = In[$signed(P[901-:32]) - 1];
			always @(*) Sgn = sv2v_tmp_CA8B4;
			wire [$signed(P[805-:32]):1] sv2v_tmp_F9BCA;
			assign sv2v_tmp_F9BCA = In[$signed(P[805-:32]) - 1:0];
			always @(*) Frac = sv2v_tmp_F9BCA;
			wire [1:1] sv2v_tmp_580D8;
			assign sv2v_tmp_580D8 = |In[$signed(P[901-:32]) - 2:$signed(P[805-:32])];
			always @(*) ExpNonZero = sv2v_tmp_580D8;
			wire [$signed(P[837-:32]):1] sv2v_tmp_2A63A;
			assign sv2v_tmp_2A63A = {In[$signed(P[901-:32]) - 2:$signed(P[805-:32]) + 1], In[$signed(P[805-:32])] | ~ExpNonZero};
			always @(*) Exp = sv2v_tmp_2A63A;
			wire [1:1] sv2v_tmp_6C177;
			assign sv2v_tmp_6C177 = &In[$signed(P[901-:32]) - 2:$signed(P[805-:32])];
			always @(*) ExpMax = sv2v_tmp_6C177;
			wire [$signed(P[901-:32]):1] sv2v_tmp_301EE;
			assign sv2v_tmp_301EE = In;
			always @(*) PostBox = sv2v_tmp_301EE;
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk1
			wire [1:1] sv2v_tmp_B03EA;
			assign sv2v_tmp_B03EA = ~(Fmt | &In[$signed(P[901-:32]) - 1:$signed(P[675-:32])]);
			always @(*) BadNaNBox = sv2v_tmp_B03EA;
			always @(*) begin
				if (_sv2v_0)
					;
				if (BadNaNBox)
					PostBox = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 1'b1, {$signed(P[643-:32]) + 1 {1'b1}}, {($signed(P[675-:32]) - $signed(P[643-:32])) - 2 {1'b0}}};
				else
					PostBox = In;
			end
			wire [1:1] sv2v_tmp_C2B86;
			assign sv2v_tmp_C2B86 = (Fmt ? In[$signed(P[901-:32]) - 1] : (BadNaNBox ? 0 : In[$signed(P[675-:32]) - 1]));
			always @(*) Sgn = sv2v_tmp_C2B86;
			wire [$signed(P[805-:32]):1] sv2v_tmp_BF14F;
			assign sv2v_tmp_BF14F = (Fmt ? In[$signed(P[805-:32]) - 1:0] : {In[$signed(P[611-:32]) - 1:0], sv2v_cast_302A5_signed(0)});
			always @(*) Frac = sv2v_tmp_BF14F;
			wire [1:1] sv2v_tmp_A4B84;
			assign sv2v_tmp_A4B84 = (Fmt ? |In[$signed(P[901-:32]) - 2:$signed(P[805-:32])] : |In[$signed(P[675-:32]) - 2:$signed(P[611-:32])]);
			always @(*) ExpNonZero = sv2v_tmp_A4B84;
			wire [$signed(P[837-:32]):1] sv2v_tmp_5869D;
			assign sv2v_tmp_5869D = (Fmt ? {In[$signed(P[901-:32]) - 2:$signed(P[805-:32]) + 1], In[$signed(P[805-:32])] | ~ExpNonZero} : {In[$signed(P[675-:32]) - 2], {$signed(P[837-:32]) - $signed(P[643-:32]) {~In[$signed(P[675-:32]) - 2]}}, In[$signed(P[675-:32]) - 3:$signed(P[611-:32]) + 1], In[$signed(P[611-:32])] | ~ExpNonZero});
			always @(*) Exp = sv2v_tmp_5869D;
			wire [1:1] sv2v_tmp_5C571;
			assign sv2v_tmp_5C571 = (Fmt ? &In[$signed(P[901-:32]) - 2:$signed(P[805-:32])] : &In[$signed(P[675-:32]) - 2:$signed(P[611-:32])]);
			always @(*) ExpMax = sv2v_tmp_5C571;
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					P[773-:2]: BadNaNBox = 1'b0;
					P[579-:2]: BadNaNBox = ~&In[$signed(P[901-:32]) - 1:$signed(P[675-:32])];
					P[449-:2]: BadNaNBox = ~&In[$signed(P[901-:32]) - 1:$signed(P[545-:32])];
					default: BadNaNBox = 1'bx;
				endcase
			end
			always @(*) begin
				if (_sv2v_0)
					;
				if (BadNaNBox & (Fmt == P[579-:2]))
					PostBox = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 1'b1, {$signed(P[643-:32]) + 1 {1'b1}}, {($signed(P[675-:32]) - $signed(P[643-:32])) - 2 {1'b0}}};
				else if (BadNaNBox)
					PostBox = {{$signed(P[901-:32]) - $signed(P[545-:32]) {1'b1}}, 1'b1, {$signed(P[513-:32]) + 1 {1'b1}}, {($signed(P[545-:32]) - $signed(P[513-:32])) - 2 {1'b0}}};
				else
					PostBox = In;
			end
			always @(*) begin
				if (_sv2v_0)
					;
				if (BadNaNBox)
					Sgn = 1'b0;
				else
					case (Fmt)
						P[773-:2]: Sgn = In[$signed(P[901-:32]) - 1];
						P[579-:2]: Sgn = In[$signed(P[675-:32]) - 1];
						P[449-:2]: Sgn = In[$signed(P[545-:32]) - 1];
						default: Sgn = 1'bx;
					endcase
			end
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					P[773-:2]: Frac = In[$signed(P[805-:32]) - 1:0];
					P[579-:2]: Frac = {In[$signed(P[611-:32]) - 1:0], sv2v_cast_302A5_signed(0)};
					P[449-:2]: Frac = {In[$signed(P[481-:32]) - 1:0], sv2v_cast_8BF36_signed(0)};
					default: Frac = {$signed(P[805-:32]) {1'bx}};
				endcase
			end
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					P[773-:2]: ExpNonZero = |In[$signed(P[901-:32]) - 2:$signed(P[805-:32])];
					P[579-:2]: ExpNonZero = |In[$signed(P[675-:32]) - 2:$signed(P[611-:32])];
					P[449-:2]: ExpNonZero = |In[$signed(P[545-:32]) - 2:$signed(P[481-:32])];
					default: ExpNonZero = 1'bx;
				endcase
			end
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					P[773-:2]: Exp = {In[$signed(P[901-:32]) - 2:$signed(P[805-:32]) + 1], In[$signed(P[805-:32])] | ~ExpNonZero};
					P[579-:2]: Exp = {In[$signed(P[675-:32]) - 2], {$signed(P[837-:32]) - $signed(P[643-:32]) {~In[$signed(P[675-:32]) - 2]}}, In[$signed(P[675-:32]) - 3:$signed(P[611-:32]) + 1], In[$signed(P[611-:32])] | ~ExpNonZero};
					P[449-:2]: Exp = {In[$signed(P[545-:32]) - 2], {$signed(P[837-:32]) - $signed(P[513-:32]) {~In[$signed(P[545-:32]) - 2]}}, In[$signed(P[545-:32]) - 3:$signed(P[481-:32]) + 1], In[$signed(P[481-:32])] | ~ExpNonZero};
					default: Exp = {$signed(P[837-:32]) {1'bx}};
				endcase
			end
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					P[773-:2]: ExpMax = &In[$signed(P[901-:32]) - 2:$signed(P[805-:32])];
					P[579-:2]: ExpMax = &In[$signed(P[675-:32]) - 2:$signed(P[611-:32])];
					P[449-:2]: ExpMax = &In[$signed(P[545-:32]) - 2:$signed(P[481-:32])];
					default: ExpMax = 1'bx;
				endcase
			end
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					2'b11: BadNaNBox = 1'b0;
					2'b01: BadNaNBox = ~&In[$signed(P[1421-:32]) - 1:$signed(P[1291-:32])];
					2'b00: BadNaNBox = ~&In[$signed(P[1421-:32]) - 1:$signed(P[1161-:32])];
					2'b10: BadNaNBox = ~&In[$signed(P[1421-:32]) - 1:$signed(P[1031-:32])];
				endcase
			end
			always @(*) begin
				if (_sv2v_0)
					;
				if (BadNaNBox)
					case (Fmt)
						2'b11: PostBox = In;
						2'b01: PostBox = {{$signed(P[1421-:32]) - $signed(P[1291-:32]) {1'b1}}, 1'b1, {$signed(P[1259-:32]) + 1 {1'b1}}, {($signed(P[1291-:32]) - $signed(P[1259-:32])) - 2 {1'b0}}};
						2'b00: PostBox = {{$signed(P[1421-:32]) - $signed(P[1161-:32]) {1'b1}}, 1'b1, {$signed(P[1129-:32]) + 1 {1'b1}}, {($signed(P[1161-:32]) - $signed(P[1129-:32])) - 2 {1'b0}}};
						2'b10: PostBox = {{$signed(P[1421-:32]) - $signed(P[1031-:32]) {1'b1}}, 1'b1, {$signed(P[999-:32]) + 1 {1'b1}}, {($signed(P[1031-:32]) - $signed(P[999-:32])) - 2 {1'b0}}};
					endcase
				else
					PostBox = In;
			end
			always @(*) begin
				if (_sv2v_0)
					;
				if (BadNaNBox)
					Sgn = 1'b0;
				else
					case (Fmt)
						2'b11: Sgn = In[$signed(P[1421-:32]) - 1];
						2'b01: Sgn = In[$signed(P[1291-:32]) - 1];
						2'b00: Sgn = In[$signed(P[1161-:32]) - 1];
						2'b10: Sgn = In[$signed(P[1031-:32]) - 1];
					endcase
			end
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					2'b11: Frac = In[$signed(P[1357-:32]) - 1:0];
					2'b01: Frac = {In[$signed(P[1227-:32]) - 1:0], sv2v_cast_FEE12_signed(0)};
					2'b00: Frac = {In[$signed(P[1097-:32]) - 1:0], sv2v_cast_E94E5_signed(0)};
					2'b10: Frac = {In[$signed(P[967-:32]) - 1:0], sv2v_cast_A7C1E_signed(0)};
				endcase
			end
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					2'b11: ExpNonZero = |In[$signed(P[1421-:32]) - 2:$signed(P[1357-:32])];
					2'b01: ExpNonZero = |In[$signed(P[1291-:32]) - 2:$signed(P[1227-:32])];
					2'b00: ExpNonZero = |In[$signed(P[1161-:32]) - 2:$signed(P[1097-:32])];
					2'b10: ExpNonZero = |In[$signed(P[1031-:32]) - 2:$signed(P[967-:32])];
				endcase
			end
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					2'b11: Exp = {In[$signed(P[1421-:32]) - 2:$signed(P[1357-:32]) + 1], In[$signed(P[1357-:32])] | ~ExpNonZero};
					2'b01: Exp = {In[$signed(P[1291-:32]) - 2], {$signed(P[1389-:32]) - $signed(P[1259-:32]) {~In[$signed(P[1291-:32]) - 2]}}, In[$signed(P[1291-:32]) - 3:$signed(P[1227-:32]) + 1], In[$signed(P[1227-:32])] | ~ExpNonZero};
					2'b00: Exp = {In[$signed(P[1161-:32]) - 2], {$signed(P[1389-:32]) - $signed(P[1129-:32]) {~In[$signed(P[1161-:32]) - 2]}}, In[$signed(P[1161-:32]) - 3:$signed(P[1097-:32]) + 1], In[$signed(P[1097-:32])] | ~ExpNonZero};
					2'b10: Exp = {In[$signed(P[1031-:32]) - 2], {$signed(P[1389-:32]) - $signed(P[999-:32]) {~In[$signed(P[1031-:32]) - 2]}}, In[$signed(P[1031-:32]) - 3:$signed(P[967-:32]) + 1], In[$signed(P[967-:32])] | ~ExpNonZero};
				endcase
			end
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					2'b11: ExpMax = &In[$signed(P[1421-:32]) - 2:$signed(P[1357-:32])];
					2'b01: ExpMax = &In[$signed(P[1291-:32]) - 2:$signed(P[1227-:32])];
					2'b00: ExpMax = &In[$signed(P[1161-:32]) - 2:$signed(P[1097-:32])];
					2'b10: ExpMax = &In[$signed(P[1031-:32]) - 2:$signed(P[967-:32])];
				endcase
			end
		end
	endgenerate
	assign FracZero = ~|Frac & ~BadNaNBox;
	assign Man = {ExpNonZero, Frac};
	assign NaN = ((ExpMax & ~FracZero) | BadNaNBox) & En;
	assign SNaN = (NaN & ~Frac[$signed(P[805-:32]) - 1]) & ~BadNaNBox;
	assign Inf = (ExpMax & FracZero) & En;
	assign Zero = ~ExpNonZero & FracZero;
	assign Subnorm = (~ExpNonZero & ~FracZero) & ~BadNaNBox;
	initial _sv2v_0 = 0;
endmodule
module adder (
	a,
	b,
	y
);
	parameter WIDTH = 8;
	input wire [WIDTH - 1:0] a;
	input wire [WIDTH - 1:0] b;
	output wire [WIDTH - 1:0] y;
	assign y = a + b;
endmodule
module aplusbeq0 (
	a,
	b,
	zero
);
	parameter WIDTH = 8;
	input wire [WIDTH - 1:0] a;
	input wire [WIDTH - 1:0] b;
	output wire zero;
	wire [WIDTH - 1:0] x;
	wire [WIDTH - 1:0] orshift;
	assign x = a ^ b;
	assign orshift = {a[WIDTH - 2:0] | b[WIDTH - 2:0], 1'b0};
	assign zero = x == orshift;
endmodule
module arrs (
	clk,
	areset,
	reset
);
	input wire clk;
	input wire areset;
	output wire reset;
	reg metaStable;
	reg resetB;
	always @(posedge clk or posedge areset)
		if (areset) begin
			metaStable <= 1'b0;
			resetB <= 1'b0;
		end
		else begin
			metaStable <= 1'b1;
			resetB <= metaStable;
		end
	assign reset = ~resetB;
endmodule
module binencoder (
	A,
	Y
);
	reg _sv2v_0;
	parameter N = 8;
	input wire [N - 1:0] A;
	output reg [$clog2(N) - 1:0] Y;
	integer index;
	always @(*) begin
		if (_sv2v_0)
			;
		Y = 1'sb0;
		for (index = 0; index < N; index = index + 1)
			if (A[index] == 1'b1)
				Y = index[$clog2(N) - 1:0];
	end
	initial _sv2v_0 = 0;
endmodule
module counter (
	clk,
	reset,
	en,
	q
);
	parameter WIDTH = 8;
	input wire clk;
	input wire reset;
	input wire en;
	output wire [WIDTH - 1:0] q;
	wire [WIDTH - 1:0] qnext;
	assign qnext = q + 1;
	flopenr #(.WIDTH(WIDTH)) cntrflop(
		.clk(clk),
		.reset(reset),
		.en(en),
		.d(qnext),
		.q(q)
	);
endmodule
module csa (
	x,
	y,
	z,
	cin,
	s,
	c
);
	parameter N = 16;
	input wire [N - 1:0] x;
	input wire [N - 1:0] y;
	input wire [N - 1:0] z;
	input wire cin;
	output wire [N - 1:0] s;
	output wire [N - 1:0] c;
	assign s = (x ^ y) ^ z;
	assign c = {(x[N - 2:0] & (y[N - 2:0] | z[N - 2:0])) | (y[N - 2:0] & z[N - 2:0]), cin};
endmodule
module decoder (
	binary,
	onehot
);
	parameter BINARY_BITS = 3;
	input wire [BINARY_BITS - 1:0] binary;
	output wire [(2 ** BINARY_BITS) - 1:0] onehot;
	assign onehot = 1 << binary;
endmodule
module mux2 (
	d0,
	d1,
	s,
	y
);
	parameter WIDTH = 8;
	input wire [WIDTH - 1:0] d0;
	input wire [WIDTH - 1:0] d1;
	input wire s;
	output wire [WIDTH - 1:0] y;
	assign y = (s ? d1 : d0);
endmodule
module mux3 (
	d0,
	d1,
	d2,
	s,
	y
);
	parameter WIDTH = 8;
	input wire [WIDTH - 1:0] d0;
	input wire [WIDTH - 1:0] d1;
	input wire [WIDTH - 1:0] d2;
	input wire [1:0] s;
	output wire [WIDTH - 1:0] y;
	assign y = (s[1] ? d2 : (s[0] ? d1 : d0));
endmodule
module mux4 (
	d0,
	d1,
	d2,
	d3,
	s,
	y
);
	parameter WIDTH = 8;
	input wire [WIDTH - 1:0] d0;
	input wire [WIDTH - 1:0] d1;
	input wire [WIDTH - 1:0] d2;
	input wire [WIDTH - 1:0] d3;
	input wire [1:0] s;
	output wire [WIDTH - 1:0] y;
	assign y = (s[1] ? (s[0] ? d3 : d2) : (s[0] ? d1 : d0));
endmodule
module mux5 (
	d0,
	d1,
	d2,
	d3,
	d4,
	s,
	y
);
	parameter WIDTH = 8;
	input wire [WIDTH - 1:0] d0;
	input wire [WIDTH - 1:0] d1;
	input wire [WIDTH - 1:0] d2;
	input wire [WIDTH - 1:0] d3;
	input wire [WIDTH - 1:0] d4;
	input wire [2:0] s;
	output wire [WIDTH - 1:0] y;
	assign y = (s[2] ? d4 : (s[1] ? (s[0] ? d3 : d2) : (s[0] ? d1 : d0)));
endmodule
module mux6 (
	d0,
	d1,
	d2,
	d3,
	d4,
	d5,
	s,
	y
);
	parameter WIDTH = 8;
	input wire [WIDTH - 1:0] d0;
	input wire [WIDTH - 1:0] d1;
	input wire [WIDTH - 1:0] d2;
	input wire [WIDTH - 1:0] d3;
	input wire [WIDTH - 1:0] d4;
	input wire [WIDTH - 1:0] d5;
	input wire [2:0] s;
	output wire [WIDTH - 1:0] y;
	assign y = (s[2] ? (s[0] ? d5 : d4) : (s[1] ? (s[0] ? d3 : d2) : (s[0] ? d1 : d0)));
endmodule
module mux7 (
	d0,
	d1,
	d2,
	d3,
	d4,
	d5,
	d6,
	s,
	y
);
	parameter WIDTH = 8;
	input wire [WIDTH - 1:0] d0;
	input wire [WIDTH - 1:0] d1;
	input wire [WIDTH - 1:0] d2;
	input wire [WIDTH - 1:0] d3;
	input wire [WIDTH - 1:0] d4;
	input wire [WIDTH - 1:0] d5;
	input wire [WIDTH - 1:0] d6;
	input wire [2:0] s;
	output wire [WIDTH - 1:0] y;
	assign y = (s[2] ? (s[1] ? d6 : (s[0] ? d5 : d4)) : (s[1] ? (s[0] ? d3 : d2) : (s[0] ? d1 : d0)));
endmodule
module neg (
	a,
	y
);
	parameter WIDTH = 8;
	input wire [WIDTH - 1:0] a;
	output wire [WIDTH - 1:0] y;
	assign y = ~a + 1;
endmodule
module onehotdecoder (
	bin,
	decoded
);
	reg _sv2v_0;
	parameter WIDTH = 2;
	input wire [WIDTH - 1:0] bin;
	output reg [(2 ** WIDTH) - 1:0] decoded;
	always @(*) begin
		if (_sv2v_0)
			;
		decoded = 1'sb0;
		decoded[bin] = 1'b1;
	end
	initial _sv2v_0 = 0;
endmodule
module or_rows (
	a,
	y
);
	parameter ROWS = 8;
	parameter COLS = 2;
	input wire [(ROWS * COLS) - 1:0] a;
	output wire [COLS - 1:0] y;
	genvar _gv_row_2;
	generate
		if (ROWS == 1) begin : genblk1
			assign y = a[0+:COLS];
		end
		else begin : genblk1
			wire [COLS - 1:0] mid [ROWS - 1:1];
			assign mid[1] = a[0+:COLS] | a[COLS+:COLS];
			for (_gv_row_2 = 2; _gv_row_2 < ROWS; _gv_row_2 = _gv_row_2 + 1) begin : genblk1
				localparam row = _gv_row_2;
				assign mid[row] = mid[row - 1] | a[row * COLS+:COLS];
			end
			assign y = mid[ROWS - 1];
		end
	endgenerate
endmodule
module priorityonehot (
	a,
	y
);
	parameter N = 8;
	input wire [N - 1:0] a;
	output wire [N - 1:0] y;
	genvar _gv_i_1;
	assign y[0] = a[0];
	generate
		for (_gv_i_1 = 1; _gv_i_1 < N; _gv_i_1 = _gv_i_1 + 1) begin : poh
			localparam i = _gv_i_1;
			assign y[i] = a[i] & ~|a[i - 1:0];
		end
	endgenerate
endmodule
module prioritythermometer (
	a,
	y
);
	parameter N = 8;
	input wire [N - 1:0] a;
	output wire [N - 1:0] y;
	genvar _gv_i_2;
	assign y[0] = ~a[0];
	generate
		for (_gv_i_2 = 1; _gv_i_2 < N; _gv_i_2 = _gv_i_2 + 1) begin : therm
			localparam i = _gv_i_2;
			assign y[i] = y[i - 1] & ~a[i];
		end
	endgenerate
endmodule
module lzc (
	num,
	ZeroCnt
);
	parameter WIDTH = 1;
	parameter CBITS = $clog2(WIDTH + 1);
	input wire [WIDTH - 1:0] num;
	output wire [CBITS - 1:0] ZeroCnt;
	wire [(WIDTH / 2) - 1:0] Lnum;
	wire [(WIDTH / 2) - 1:0] Rnum;
	wire [CBITS - 2:0] LCnt;
	wire [CBITS - 2:0] RCnt;
	assign Lnum = num[WIDTH - 1-:WIDTH / 2];
	assign Rnum = num[(WIDTH / 2) - 1-:WIDTH / 2];
	generate
		if (WIDTH <= 2) begin : genblk1
			assign ZeroCnt = (num == 2'b00 ? 2'b10 : (num == 2'b01 ? 2'b01 : 2'b00));
		end
		else begin : genblk1
			lzc #(.WIDTH(WIDTH / 2)) l_lcz(
				.num(Lnum),
				.ZeroCnt(LCnt)
			);
			lzc #(.WIDTH(WIDTH / 2)) r_lcz(
				.num(Rnum),
				.ZeroCnt(RCnt)
			);
			assign ZeroCnt = (~LCnt[CBITS - 2] ? {LCnt[CBITS - 2] & RCnt[CBITS - 2], 1'b0, LCnt[CBITS - 3:0]} : {LCnt[CBITS - 2] & RCnt[CBITS - 2], ~RCnt[CBITS - 2], RCnt[CBITS - 3:0]});
		end
	endgenerate
endmodule
module hazard (
	BPWrongE,
	CSRWriteFenceM,
	RetM,
	TrapM,
	StructuralStallD,
	LSUStallM,
	IFUStallF,
	FPUStallD,
	ExternalStall,
	DivBusyE,
	FDivBusyE,
	wfiM,
	IntPendingM,
	StallF,
	StallD,
	StallE,
	StallM,
	StallW,
	FlushD,
	FlushE,
	FlushM,
	FlushW
);
	input wire BPWrongE;
	input wire CSRWriteFenceM;
	input wire RetM;
	input wire TrapM;
	input wire StructuralStallD;
	input wire LSUStallM;
	input wire IFUStallF;
	input wire FPUStallD;
	input wire ExternalStall;
	input wire DivBusyE;
	input wire FDivBusyE;
	input wire wfiM;
	input wire IntPendingM;
	output wire StallF;
	output wire StallD;
	output wire StallE;
	output wire StallM;
	output wire StallW;
	output wire FlushD;
	output wire FlushE;
	output wire FlushM;
	output wire FlushW;
	wire StallFCause;
	wire StallDCause;
	wire StallECause;
	wire StallMCause;
	wire StallWCause;
	wire LatestUnstalledD;
	wire LatestUnstalledE;
	wire LatestUnstalledM;
	wire LatestUnstalledW;
	wire FlushDCause;
	wire FlushECause;
	wire FlushMCause;
	wire FlushWCause;
	wire WFIStallM;
	wire WFIInterruptedM;
	assign WFIStallM = wfiM & ~IntPendingM;
	assign WFIInterruptedM = wfiM & IntPendingM;
	assign FlushDCause = ((TrapM | RetM) | CSRWriteFenceM) | BPWrongE;
	assign FlushECause = ((TrapM | RetM) | CSRWriteFenceM) | (BPWrongE & ~(DivBusyE | FDivBusyE));
	assign FlushMCause = (TrapM | RetM) | CSRWriteFenceM;
	assign FlushWCause = TrapM & ~WFIInterruptedM;
	assign StallFCause = 1'b0;
	assign StallDCause = (StructuralStallD | FPUStallD) & ~FlushDCause;
	assign StallECause = (DivBusyE | FDivBusyE) & ~FlushECause;
	assign StallMCause = WFIStallM & ~FlushMCause;
	assign StallWCause = ((IFUStallF & ~FlushDCause) | (LSUStallM & ~FlushWCause)) | ExternalStall;
	assign StallF = StallFCause | StallD;
	assign StallD = StallDCause | StallE;
	assign StallE = StallECause | StallM;
	assign StallM = StallMCause | StallW;
	assign StallW = StallWCause;
	assign LatestUnstalledD = ~StallD & StallF;
	assign LatestUnstalledE = ~StallE & StallD;
	assign LatestUnstalledM = ~StallM & StallE;
	assign LatestUnstalledW = ~StallW & StallM;
	assign FlushD = LatestUnstalledD | FlushDCause;
	assign FlushE = LatestUnstalledE | FlushECause;
	assign FlushM = LatestUnstalledM | FlushMCause;
	assign FlushW = LatestUnstalledW | FlushWCause;
endmodule
module alu (
	A,
	B,
	W64,
	UW64,
	SubArith,
	ALUSelect,
	BSelect,
	ZBBSelect,
	Funct3,
	Funct7,
	Rs2E,
	BALUControl,
	BMUActive,
	CZero,
	ALUResult,
	Sum
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[4216-:32]) - 1:0] A;
	input wire [$signed(P[4216-:32]) - 1:0] B;
	input wire W64;
	input wire UW64;
	input wire SubArith;
	input wire [2:0] ALUSelect;
	input wire [3:0] BSelect;
	input wire [3:0] ZBBSelect;
	input wire [2:0] Funct3;
	input wire [6:0] Funct7;
	input wire [4:0] Rs2E;
	input wire [2:0] BALUControl;
	input wire BMUActive;
	input wire [1:0] CZero;
	output wire [$signed(P[4216-:32]) - 1:0] ALUResult;
	output wire [$signed(P[4216-:32]) - 1:0] Sum;
	wire [$signed(P[4216-:32]) - 1:0] CondMaskInvB;
	wire [$signed(P[4216-:32]) - 1:0] Shift;
	reg [$signed(P[4216-:32]) - 1:0] FullResult;
	wire [$signed(P[4216-:32]) - 1:0] PreALUResult;
	wire [$signed(P[4216-:32]) - 1:0] CondMaskB;
	wire [$signed(P[4216-:32]) - 1:0] CondShiftA;
	reg [$signed(P[4216-:32]) - 1:0] ZeroCondMaskInvB;
	wire [$signed(P[4216-:32]) - 1:0] AndResult;
	wire Carry;
	wire Neg;
	wire LT;
	wire LTU;
	wire Asign;
	wire Bsign;
	assign CondMaskInvB = (SubArith ? ~CondMaskB : CondMaskB);
	assign {Carry, Sum} = (CondShiftA + CondMaskInvB) + {{$signed(P[4216-:32]) - 1 {1'b0}}, SubArith};
	generate
		if (P[4058]) begin : zicond
			wire BZero;
			assign BZero = B == 0;
			always @(*) begin
				if (_sv2v_0)
					;
				case (CZero)
					2'b01: ZeroCondMaskInvB = {$signed(P[4216-:32]) {~BZero}};
					2'b10: ZeroCondMaskInvB = {$signed(P[4216-:32]) {BZero}};
					default: ZeroCondMaskInvB = CondMaskInvB;
				endcase
			end
		end
		else begin : genblk1
			wire [$signed(P[4216-:32]):1] sv2v_tmp_C8935;
			assign sv2v_tmp_C8935 = CondMaskInvB;
			always @(*) ZeroCondMaskInvB = sv2v_tmp_C8935;
		end
	endgenerate
	shifter #(.P(P)) sh(
		.A(CondShiftA),
		.Amt(B[$signed(P[1485-:32]) - 1:0]),
		.Right(Funct3[2]),
		.W64(W64),
		.SubArith(SubArith),
		.Y(Shift),
		.Rotate(BALUControl[2])
	);
	assign Neg = Sum[$signed(P[4216-:32]) - 1];
	assign Asign = A[$signed(P[4216-:32]) - 1];
	assign Bsign = B[$signed(P[4216-:32]) - 1];
	assign LT = ((Asign & ~Bsign) | (Asign & Neg)) | (~Bsign & Neg);
	assign LTU = ~Carry;
	assign AndResult = A & ZeroCondMaskInvB;
	always @(*) begin
		if (_sv2v_0)
			;
		case (ALUSelect)
			3'b000: FullResult = Sum;
			3'b001: FullResult = Shift;
			3'b010: FullResult = {{$signed(P[4216-:32]) - 1 {1'b0}}, LT};
			3'b011: FullResult = {{$signed(P[4216-:32]) - 1 {1'b0}}, LTU};
			3'b100: FullResult = A ^ CondMaskInvB;
			3'b101: FullResult = (P[1755] ? {{$signed(P[4216-:32]) - 1 {1'b0}}, |AndResult} : Shift);
			3'b110: FullResult = A | CondMaskInvB;
			3'b111: FullResult = AndResult;
		endcase
	end
	generate
		if ($signed(P[4216-:32]) == 64) begin : genblk2
			assign PreALUResult = (W64 ? {{32 {FullResult[31]}}, FullResult[31:0]} : FullResult);
		end
		else begin : genblk2
			assign PreALUResult = FullResult;
		end
		if (((((((((P[1756] | P[1755]) | P[1758]) | P[1757]) | P[1750]) | P[1749]) | P[1748]) | P[1747]) | P[1746]) | P[1745]) begin : bitmanipalu
			bitmanipalu #(.P(P)) balu(
				.A(A),
				.B(B),
				.W64(W64),
				.UW64(UW64),
				.BSelect(BSelect),
				.ZBBSelect(ZBBSelect),
				.BMUActive(BMUActive),
				.Funct3(Funct3),
				.Funct7(Funct7),
				.Rs2E(Rs2E),
				.LT(LT),
				.LTU(LTU),
				.BALUControl(BALUControl),
				.PreALUResult(PreALUResult),
				.FullResult(FullResult),
				.CondMaskB(CondMaskB),
				.CondShiftA(CondShiftA),
				.ALUResult(ALUResult)
			);
		end
		else begin : genblk3
			assign ALUResult = PreALUResult;
			assign CondMaskB = B;
			assign CondShiftA = A;
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module comparator (
	a,
	b,
	sgnd,
	flags
);
	parameter WIDTH = 64;
	input wire [WIDTH - 1:0] a;
	input wire [WIDTH - 1:0] b;
	input wire sgnd;
	output wire [1:0] flags;
	wire eq;
	wire lt;
	wire [WIDTH - 1:0] af;
	wire [WIDTH - 1:0] bf;
	assign af = {a[WIDTH - 1] ^ sgnd, a[WIDTH - 2:0]};
	assign bf = {b[WIDTH - 1] ^ sgnd, b[WIDTH - 2:0]};
	assign eq = a == b;
	assign lt = af < bf;
	assign flags = {eq, lt};
endmodule
module controller (
	clk,
	reset,
	StallD,
	FlushD,
	InstrD,
	STATUS_FS,
	ENVCFG_CBE,
	ImmSrcD,
	IllegalIEUFPUInstrD,
	IllegalBaseInstrD,
	JumpD,
	BranchD,
	StructuralStallD,
	LoadStallD,
	StoreStallD,
	Rs1D,
	Rs2D,
	Rs2E,
	StallE,
	FlushE,
	FlagsE,
	FWriteIntE,
	FCvtIntE,
	PCSrcE,
	ALUSrcAE,
	ALUSrcBE,
	ALUResultSrcE,
	ALUSelectE,
	Funct3E,
	Funct7E,
	IntDivE,
	W64E,
	UW64E,
	SubArithE,
	JumpE,
	BranchE,
	BranchSignedE,
	BSelectE,
	ZBBSelectE,
	BALUControlE,
	BMUActiveE,
	CZeroE,
	MDUActiveE,
	CMOpM,
	IFUPrefetchE,
	LSUPrefetchM,
	ForwardAE,
	ForwardBE,
	StallM,
	FlushM,
	MemRWE,
	MemRWM,
	CSRReadM,
	CSRWriteM,
	PrivilegedM,
	AtomicM,
	Funct3M,
	InvalidateICacheM,
	FlushDCacheM,
	InstrValidD,
	InstrValidE,
	InstrValidM,
	FWriteIntM,
	StallW,
	FlushW,
	RegWriteW,
	IntDivW,
	ResultSrcW,
	CSRWriteFenceM,
	RdE,
	RdM,
	RdW
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallD;
	input wire FlushD;
	input wire [31:0] InstrD;
	input wire [1:0] STATUS_FS;
	input wire [3:0] ENVCFG_CBE;
	output reg [2:0] ImmSrcD;
	input wire IllegalIEUFPUInstrD;
	output wire IllegalBaseInstrD;
	output wire JumpD;
	output wire BranchD;
	output wire StructuralStallD;
	output wire LoadStallD;
	output wire StoreStallD;
	output wire [4:0] Rs1D;
	output wire [4:0] Rs2D;
	output wire [4:0] Rs2E;
	input wire StallE;
	input wire FlushE;
	input wire [1:0] FlagsE;
	input wire FWriteIntE;
	input wire FCvtIntE;
	output wire PCSrcE;
	output wire ALUSrcAE;
	output wire ALUSrcBE;
	output wire ALUResultSrcE;
	output wire [2:0] ALUSelectE;
	output wire [2:0] Funct3E;
	output wire [6:0] Funct7E;
	output wire IntDivE;
	output wire W64E;
	output wire UW64E;
	output wire SubArithE;
	output wire JumpE;
	output wire BranchE;
	output wire BranchSignedE;
	output wire [3:0] BSelectE;
	output wire [3:0] ZBBSelectE;
	output wire [2:0] BALUControlE;
	output wire BMUActiveE;
	output wire [1:0] CZeroE;
	output wire MDUActiveE;
	output wire [3:0] CMOpM;
	output wire IFUPrefetchE;
	output wire LSUPrefetchM;
	output reg [1:0] ForwardAE;
	output reg [1:0] ForwardBE;
	input wire StallM;
	input wire FlushM;
	output wire [1:0] MemRWE;
	output wire [1:0] MemRWM;
	output wire CSRReadM;
	output wire CSRWriteM;
	output wire PrivilegedM;
	output wire [1:0] AtomicM;
	output wire [2:0] Funct3M;
	output wire InvalidateICacheM;
	output wire FlushDCacheM;
	output wire InstrValidD;
	output wire InstrValidE;
	output wire InstrValidM;
	output wire FWriteIntM;
	input wire StallW;
	input wire FlushW;
	output wire RegWriteW;
	output wire IntDivW;
	output wire [2:0] ResultSrcW;
	output wire CSRWriteFenceM;
	output wire [4:0] RdE;
	output wire [4:0] RdM;
	output wire [4:0] RdW;
	wire [4:0] Rs1E;
	wire [6:0] OpD;
	wire [2:0] Funct3D;
	wire [6:0] Funct7D;
	wire [4:0] RdD;
	wire RegWriteD;
	wire RegWriteE;
	wire [2:0] ResultSrcD;
	wire [2:0] ResultSrcE;
	wire [2:0] ResultSrcM;
	wire [2:0] PreImmSrcD;
	wire [1:0] MemRWD;
	wire ALUOpD;
	wire BaseW64D;
	wire BaseRegWriteD;
	wire BaseSubArithD;
	wire BaseALUSrcBD;
	wire ALUSrcAD;
	wire ALUSrcBD;
	wire ALUResultSrcD;
	wire W64D;
	wire MDUD;
	wire CSRZeroSrcD;
	wire CSRReadD;
	wire [1:0] AtomicD;
	wire FenceXD;
	wire CMOD;
	wire InvalidateICacheD;
	wire FlushDCacheD;
	wire MemReadE;
	wire CSRReadE;
	wire MDUE;
	wire SCE;
	wire CSRWriteD;
	wire CSRWriteE;
	wire PrivilegedD;
	wire PrivilegedE;
	wire InvalidateICacheE;
	wire FlushDCacheE;
	reg [23:0] ControlsD;
	wire SubArithD;
	wire subD;
	wire sraD;
	wire sltD;
	wire sltuD;
	wire BranchTakenE;
	wire eqE;
	wire ltE;
	wire unused;
	wire BranchFlagE;
	wire IEURegWriteE;
	wire IllegalERegAdrD;
	wire [1:0] AtomicE;
	wire FenceD;
	wire FenceE;
	wire SFenceVmaD;
	wire IntDivM;
	wire RegWriteM;
	wire [1:0] CZeroD;
	wire IFunctD;
	wire RFunctD;
	wire MFunctD;
	wire LFunctD;
	wire SFunctD;
	wire BFunctD;
	wire FLSFunctD;
	wire JRFunctD;
	wire FenceFunctD;
	wire CMOFunctD;
	wire AFunctD;
	wire AMOFunctD;
	wire RWFunctD;
	wire MWFunctD;
	wire PFunctD;
	wire CSRFunctD;
	wire FenceM;
	wire [2:0] PreALUSelectD;
	wire [2:0] ALUSelectD;
	wire IWValidFunct3D;
	reg [3:0] CMOpD;
	wire [3:0] CMOpE;
	reg IFUPrefetchD;
	reg LSUPrefetchD;
	wire LSUPrefetchE;
	wire MatchDE;
	wire FCvtIntStallD;
	wire MDUStallD;
	wire CSRRdStallD;
	wire FunctCZeroD;
	wire BUW64D;
	assign OpD = InstrD[6:0];
	assign Funct3D = InstrD[14:12];
	assign Funct7D = InstrD[31:25];
	assign Rs1D = InstrD[19:15];
	assign Rs2D = InstrD[24:20];
	assign RdD = InstrD[11:7];
	generate
		if (((((((((((P[4086] | P[1758]) | P[1757]) | P[1756]) | P[1755]) | P[1750]) | P[1749]) | P[1748]) | P[1746]) | P[1747]) | P[1745]) | P[4058]) begin : legalcheck
			wire Funct7ZeroD;
			wire Funct7b5D;
			wire IShiftD;
			wire INoShiftD;
			wire Funct7ShiftZeroD;
			wire Funct7Shiftb5D;
			assign Funct7ZeroD = Funct7D == 7'b0000000;
			assign Funct7b5D = Funct7D == 7'b0100000;
			assign FunctCZeroD = (((Funct3D == 3'b101) | (Funct3D == 3'b111)) & (Funct7D == 7'b0000111)) & P[4058];
			assign Funct7ShiftZeroD = (($signed(P[4216-:32]) == 64) & ~OpD[3] ? Funct7D[6:1] == 6'b000000 : Funct7ZeroD);
			assign Funct7Shiftb5D = (($signed(P[4216-:32]) == 64) & ~OpD[3] ? Funct7D[6:1] == 6'b010000 : Funct7b5D);
			assign IShiftD = ((Funct3D == 3'b001) & Funct7ShiftZeroD) | ((Funct3D == 3'b101) & (Funct7ShiftZeroD | Funct7Shiftb5D));
			assign INoShiftD = (Funct3D != 3'b001) & (Funct3D != 3'b101);
			assign IFunctD = IShiftD | INoShiftD;
			assign RFunctD = ((((Funct3D == 3'b000) | (Funct3D == 3'b101)) & Funct7b5D) | FunctCZeroD) | Funct7ZeroD;
			assign MFunctD = (Funct7D == 7'b0000001) & (P[1489] | (P[4063] & ~Funct3D[2]));
			assign LFunctD = (((((Funct3D == 3'b000) | (Funct3D == 3'b001)) | (Funct3D == 3'b010)) | (Funct3D == 3'b100)) | (Funct3D == 3'b101)) | (($signed(P[4216-:32]) == 64) & ((Funct3D == 3'b011) | (Funct3D == 3'b110)));
			assign FLSFunctD = (STATUS_FS != 2'b00) & (((((Funct3D == 3'b010) & P[1491]) | ((Funct3D == 3'b011) & P[1493])) | ((Funct3D == 3'b100) & P[1488])) | ((Funct3D == 3'b001) & P[4070]));
			assign FenceFunctD = (Funct3D == 3'b000) | (P[4085] & (Funct3D == 3'b001));
			assign CMOFunctD = ((Funct3D == 3'b010) & (RdD == 5'b00000)) & (((P[4061] & (InstrD[31:20] == 12'd4)) & ENVCFG_CBE[3]) | ((P[4062] & ((InstrD[31:20] == 12'd0) & (ENVCFG_CBE[1:0] != 2'b00))) | (((InstrD[31:20] == 12'd1) | (InstrD[31:20] == 12'd2)) & ENVCFG_CBE[2])));
			assign AFunctD = (Funct3D == 3'b010) | (($signed(P[4216-:32]) == 64) & (Funct3D == 3'b011));
			assign AMOFunctD = ((((((((InstrD[31:27] == 5'b00001) | (InstrD[31:27] == 5'b00000)) | (InstrD[31:27] == 5'b00100)) | (InstrD[31:27] == 5'b01100)) | (InstrD[31:27] == 5'b01000)) | (InstrD[31:27] == 5'b10000)) | (InstrD[31:27] == 5'b10100)) | (InstrD[31:27] == 5'b11000)) | (InstrD[31:27] == 5'b11100);
			assign RWFunctD = (((((Funct3D == 3'b000) | (Funct3D == 3'b001)) | (Funct3D == 3'b101)) & Funct7ZeroD) | (((Funct3D == 3'b000) | (Funct3D == 3'b101)) & Funct7b5D)) & ($signed(P[4216-:32]) == 64);
			assign MWFunctD = (MFunctD & ($signed(P[4216-:32]) == 64)) & ~(((Funct3D == 3'b001) | (Funct3D == 3'b010)) | (Funct3D == 3'b011));
			assign SFunctD = (((Funct3D == 3'b000) | (Funct3D == 3'b001)) | (Funct3D == 3'b010)) | (($signed(P[4216-:32]) == 64) & (Funct3D == 3'b011));
			assign BFunctD = Funct3D[2:1] != 2'b01;
			assign JRFunctD = Funct3D == 3'b000;
			assign PFunctD = (Funct3D == 3'b000) & (RdD == 5'b00000);
			assign CSRFunctD = Funct3D[1:0] != 2'b00;
			assign IWValidFunct3D = ((Funct3D == 3'b000) | (Funct3D == 3'b001)) | (Funct3D == 3'b101);
		end
		else begin : legalcheck2
			assign IFunctD = 1'b1;
			assign RFunctD = ~Funct7D[0];
			assign MFunctD = Funct7D[0] & (P[1489] | (P[4063] & ~Funct3D[2]));
			assign LFunctD = 1'b1;
			assign FLSFunctD = 1'b1;
			assign FenceFunctD = 1'b1;
			assign CMOFunctD = 1'b1;
			assign AFunctD = 1'b1;
			assign AMOFunctD = 1'b1;
			assign RWFunctD = 1'b1;
			assign MWFunctD = 1'b1;
			assign SFunctD = 1'b1;
			assign BFunctD = 1'b1;
			assign JRFunctD = 1'b1;
			assign PFunctD = 1'b1;
			assign CSRFunctD = 1'b1;
			assign IWValidFunct3D = 1'b1;
		end
	endgenerate
	always @(*) begin
		if (_sv2v_0)
			;
		ControlsD = 24'b000000000000000000000001;
		case (OpD)
			7'b0000011:
				if (LFunctD)
					ControlsD = 24'b100001100010000000000000;
			7'b0000111:
				if (FLSFunctD)
					ControlsD = 24'b000001100010000000000001;
			7'b0001111:
				if (FenceFunctD) begin
					if (P[4085])
						ControlsD = 24'b000000000000000000100000;
					else
						ControlsD = 24'b000000000000000000000000;
				end
				else if (CMOFunctD)
					ControlsD = 24'b010101000000000000000010;
			7'b0010011:
				if (IFunctD)
					ControlsD = 24'b100001000000100000000000;
			7'b0010111: ControlsD = 24'b110011000000000000000000;
			7'b0011011:
				if ((IFunctD & IWValidFunct3D) & ($signed(P[4216-:32]) == 64))
					ControlsD = 24'b100001000000100100000000;
			7'b0100011:
				if (SFunctD)
					ControlsD = 24'b000101010000000000000000;
			7'b0100111:
				if (FLSFunctD)
					ControlsD = 24'b000101010000000000000001;
			7'b0101111:
				if (AFunctD) begin
					if ((P[4053] & (InstrD[31:27] == 5'b00010)) & (Rs2D == 5'b00000))
						ControlsD = 24'b100000100010000000000100;
					else if (P[4053] & (InstrD[31:27] == 5'b00011))
						ControlsD = 24'b110101011000000000000100;
					else if (P[4054] & AMOFunctD)
						ControlsD = 24'b110101110010000000001000;
				end
			7'b0110011:
				if (RFunctD)
					ControlsD = 24'b100000000000100000000000;
				else if (MFunctD)
					ControlsD = 24'b100000000110000000010000;
			7'b0110111: ControlsD = 24'b110001000000001000000000;
			7'b0111011:
				if (RWFunctD)
					ControlsD = 24'b100000000000100100000000;
				else if (MWFunctD)
					ControlsD = 24'b100000000110000100010000;
			7'b1100011:
				if (BFunctD)
					ControlsD = 24'b001011000001000000000000;
			7'b1100111:
				if (JRFunctD)
					ControlsD = 24'b100001000000011000000000;
			7'b1101111: ControlsD = 24'b101111000000011000000000;
			7'b1110011:
				if (P[4086]) begin
					if (PFunctD)
						ControlsD = 24'b000000000000000001000000;
					else if (CSRFunctD)
						ControlsD = 24'b100000000100000010000000;
				end
		endcase
	end
	assign IllegalERegAdrD = ((P[1492] & P[4086]) & ControlsD[23]) & InstrD[11];
	assign {BaseRegWriteD, PreImmSrcD, ALUSrcAD, BaseALUSrcBD, MemRWD, ResultSrcD, BranchD, ALUOpD, JumpD, ALUResultSrcD, BaseW64D, CSRReadD, PrivilegedD, FenceXD, MDUD, AtomicD, CMOD, unused} = (IllegalIEUFPUInstrD ? 24'b000000000000000000000000 : ControlsD);
	assign CSRZeroSrcD = (InstrD[14] ? InstrD[19:15] == 0 : Rs1D == 0);
	assign CSRWriteD = CSRReadD & !(CSRZeroSrcD & InstrD[13]);
	assign SFenceVmaD = PrivilegedD & (InstrD[31:25] == 7'b0001001);
	assign FenceD = SFenceVmaD | FenceXD;
	assign sltuD = Funct3D == 3'b011;
	assign subD = ((Funct3D == 3'b000) & Funct7D[5]) & OpD[5];
	assign sraD = (Funct3D == 3'b101) & Funct7D[5];
	assign BaseSubArithD = ALUOpD & (((subD | sraD) | sltD) | sltuD);
	generate
		if (((((((((P[1755] | P[1758]) | P[1757]) | P[1756]) | P[1750]) | P[1749]) | P[1748]) | P[1746]) | P[1747]) | P[1745]) begin : bitmanipi
			wire IllegalBitmanipInstrD;
			wire BRegWriteD;
			wire BW64D;
			wire BSubArithD;
			wire BALUSrcBD;
			bmuctrl #(.P(P)) bmuctrl(
				.clk(clk),
				.reset(reset),
				.InstrD(InstrD),
				.ALUOpD(ALUOpD),
				.BRegWriteD(BRegWriteD),
				.BALUSrcBD(BALUSrcBD),
				.BW64D(BW64D),
				.BUW64D(BUW64D),
				.BSubArithD(BSubArithD),
				.IllegalBitmanipInstrD(IllegalBitmanipInstrD),
				.StallE(StallE),
				.FlushE(FlushE),
				.ALUSelectD(PreALUSelectD),
				.BSelectE(BSelectE),
				.ZBBSelectE(ZBBSelectE),
				.BALUControlE(BALUControlE),
				.BMUActiveE(BMUActiveE)
			);
			if (P[1758]) begin : genblk1
				assign sltD = (Funct3D == 3'b010) & (~Funct7D[4] | ~OpD[5]);
			end
			else begin : genblk1
				assign sltD = Funct3D == 3'b010;
			end
			assign IllegalBaseInstrD = (ControlsD[0] & IllegalBitmanipInstrD) | IllegalERegAdrD;
			assign RegWriteD = BaseRegWriteD | BRegWriteD;
			assign W64D = BaseW64D | BW64D;
			assign ALUSrcBD = BaseALUSrcBD | BALUSrcBD;
			assign SubArithD = BaseSubArithD | BSubArithD;
		end
		else begin : bitmanipi
			assign PreALUSelectD = (ALUOpD ? Funct3D : 3'b000);
			assign sltD = Funct3D == 3'b010;
			assign IllegalBaseInstrD = ControlsD[0] | IllegalERegAdrD;
			assign RegWriteD = BaseRegWriteD;
			assign W64D = BaseW64D;
			assign ALUSrcBD = BaseALUSrcBD;
			assign SubArithD = BaseSubArithD;
			assign BUW64D = 1'b0;
			assign BSelectE = 4'b0000;
			assign ZBBSelectE = 4'b0000;
			assign BALUControlE = 3'b000;
			assign BMUActiveE = 1'b0;
		end
		if (P[4058]) begin : Zicond
			wire SomeCZeroD;
			assign SomeCZeroD = FunctCZeroD & (OpD == 7'b0110011);
			assign CZeroD = {SomeCZeroD & (Funct3D == 3'b111), SomeCZeroD & (Funct3D == 3'b101)};
			assign ALUSelectD = (SomeCZeroD ? 3'b111 : PreALUSelectD);
		end
		else begin : genblk3
			assign CZeroD = 2'b00;
			assign ALUSelectD = PreALUSelectD;
		end
		if (P[4085] & (P[4050] | P[4051])) begin : fencei
			wire FenceID;
			assign FenceID = FenceXD & (Funct3D == 3'b001);
			assign InvalidateICacheD = FenceID;
			assign FlushDCacheD = FenceID;
		end
		else begin : fencei
			assign InvalidateICacheD = 1'b0;
			assign FlushDCacheD = 1'b0;
		end
	endgenerate
	always @(*) begin
		if (_sv2v_0)
			;
		CMOpD = 4'b0000;
		if (P[4061] & CMOD)
			CMOpD[3] = InstrD[31:20] == 12'd4;
		if (P[4062] & CMOD) begin
			CMOpD[2] = InstrD[31:20] == 12'd2;
			CMOpD[1] = (InstrD[31:20] == 12'd1) | ((InstrD[31:20] == 12'd0) & (ENVCFG_CBE[1:0] == 2'b01));
			CMOpD[0] = (InstrD[31:20] == 12'd0) & (ENVCFG_CBE[1:0] == 2'b11);
		end
	end
	always @(*) begin
		if (_sv2v_0)
			;
		IFUPrefetchD = 1'b0;
		LSUPrefetchD = 1'b0;
		ImmSrcD = PreImmSrcD;
		if (P[4060] & (InstrD[14:0] == 15'b110000000010011)) begin
			case (Rs2D)
				5'b00000: IFUPrefetchD = 1'b1;
				5'b00001: LSUPrefetchD = 1'b1;
				5'b00011: LSUPrefetchD = 1'b1;
			endcase
			if (IFUPrefetchD | LSUPrefetchD)
				ImmSrcD = 3'b001;
		end
	end
	flopenrc #(.WIDTH(1)) controlregD(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallD),
		.d(1'b1),
		.q(InstrValidD)
	);
	flopenrc #(.WIDTH(45)) controlregE(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d({ALUSelectD, RegWriteD, ResultSrcD, MemRWD, JumpD, BranchD, ALUSrcAD, ALUSrcBD, ALUResultSrcD, CSRReadD, CSRWriteD, PrivilegedD, Funct3D, Funct7D, W64D, BUW64D, SubArithD, MDUD, AtomicD, InvalidateICacheD, FlushDCacheD, FenceD, CMOpD, IFUPrefetchD, LSUPrefetchD, CZeroD, InstrValidD}),
		.q({ALUSelectE, IEURegWriteE, ResultSrcE, MemRWE, JumpE, BranchE, ALUSrcAE, ALUSrcBE, ALUResultSrcE, CSRReadE, CSRWriteE, PrivilegedE, Funct3E, Funct7E, W64E, UW64E, SubArithE, MDUE, AtomicE, InvalidateICacheE, FlushDCacheE, FenceE, CMOpE, IFUPrefetchE, LSUPrefetchE, CZeroE, InstrValidE})
	);
	flopenrc #(.WIDTH(5)) Rs1EReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(Rs1D),
		.q(Rs1E)
	);
	flopenrc #(.WIDTH(5)) Rs2EReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(Rs2D),
		.q(Rs2E)
	);
	flopenrc #(.WIDTH(5)) RdEReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(RdD),
		.q(RdE)
	);
	assign BranchSignedE = ~(Funct3E[2:1] == 2'b11) & BranchE;
	assign {eqE, ltE} = FlagsE;
	mux2 #(.WIDTH(1)) branchflagmux(
		.d0(eqE),
		.d1(ltE),
		.s(Funct3E[2]),
		.y(BranchFlagE)
	);
	assign BranchTakenE = BranchFlagE ^ Funct3E[0];
	assign PCSrcE = JumpE | (BranchE & BranchTakenE);
	assign MemReadE = MemRWE[1];
	assign SCE = ResultSrcE == 3'b100;
	assign MDUActiveE = ResultSrcE == 3'b011;
	assign RegWriteE = IEURegWriteE | FWriteIntE;
	assign IntDivE = MDUE & Funct3E[2];
	flopenrc #(.WIDTH(25)) controlregM(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d({RegWriteE, ResultSrcE, MemRWE, CSRReadE, CSRWriteE, PrivilegedE, Funct3E, FWriteIntE, AtomicE, InvalidateICacheE, FlushDCacheE, FenceE, InstrValidE, IntDivE, CMOpE, LSUPrefetchE}),
		.q({RegWriteM, ResultSrcM, MemRWM, CSRReadM, CSRWriteM, PrivilegedM, Funct3M, FWriteIntM, AtomicM, InvalidateICacheM, FlushDCacheM, FenceM, InstrValidM, IntDivM, CMOpM, LSUPrefetchM})
	);
	flopenrc #(.WIDTH(5)) RdMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(RdE),
		.q(RdM)
	);
	flopenrc #(.WIDTH(5)) controlregW(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d({RegWriteM, ResultSrcM, IntDivM}),
		.q({RegWriteW, ResultSrcW, IntDivW})
	);
	flopenrc #(.WIDTH(5)) RdWReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(RdM),
		.q(RdW)
	);
	assign CSRWriteFenceM = CSRWriteM | FenceM;
	always @(*) begin
		if (_sv2v_0)
			;
		ForwardAE = 2'b00;
		ForwardBE = 2'b00;
		if (Rs1E != 5'b00000) begin
			if ((Rs1E == RdM) & RegWriteM)
				ForwardAE = 2'b10;
			else if ((Rs1E == RdW) & RegWriteW)
				ForwardAE = 2'b01;
		end
		if (Rs2E != 5'b00000) begin
			if ((Rs2E == RdM) & RegWriteM)
				ForwardBE = 2'b10;
			else if ((Rs2E == RdW) & RegWriteW)
				ForwardBE = 2'b01;
		end
	end
	assign MatchDE = ((Rs1D == RdE) | (Rs2D == RdE)) & (RdE != 5'b00000);
	assign LoadStallD = (MemReadE | SCE) & MatchDE;
	assign StoreStallD = MemRWD[1] & MemRWE[0];
	assign CSRRdStallD = CSRReadE & MatchDE;
	assign MDUStallD = MDUE & MatchDE;
	assign FCvtIntStallD = FCvtIntE & MatchDE;
	assign StructuralStallD = (((LoadStallD | StoreStallD) | CSRRdStallD) | MDUStallD) | FCvtIntStallD;
	initial _sv2v_0 = 0;
endmodule
module datapath (
	clk,
	reset,
	ImmSrcD,
	InstrD,
	Rs1D,
	Rs2D,
	Rs2E,
	PCE,
	PCLinkE,
	Funct3E,
	Funct7E,
	StallE,
	FlushE,
	ForwardAE,
	ForwardBE,
	W64E,
	UW64E,
	SubArithE,
	ALUSrcAE,
	ALUSrcBE,
	ALUResultSrcE,
	ALUSelectE,
	JumpE,
	BranchSignedE,
	BSelectE,
	ZBBSelectE,
	BALUControlE,
	BMUActiveE,
	CZeroE,
	FlagsE,
	IEUAdrE,
	ForwardedSrcAE,
	ForwardedSrcBE,
	StallM,
	FlushM,
	FWriteIntM,
	FCvtIntW,
	FIntResM,
	SrcAM,
	WriteDataM,
	StallW,
	FlushW,
	RegWriteW,
	IntDivW,
	SquashSCW,
	ResultSrcW,
	FCvtIntResW,
	ReadDataW,
	CSRReadValW,
	MDUResultW,
	FIntDivResultW,
	RdW
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire [2:0] ImmSrcD;
	input wire [31:0] InstrD;
	input wire [4:0] Rs1D;
	input wire [4:0] Rs2D;
	input wire [4:0] Rs2E;
	input wire [$signed(P[4216-:32]) - 1:0] PCE;
	input wire [$signed(P[4216-:32]) - 1:0] PCLinkE;
	input wire [2:0] Funct3E;
	input wire [6:0] Funct7E;
	input wire StallE;
	input wire FlushE;
	input wire [1:0] ForwardAE;
	input wire [1:0] ForwardBE;
	input wire W64E;
	input wire UW64E;
	input wire SubArithE;
	input wire ALUSrcAE;
	input wire ALUSrcBE;
	input wire ALUResultSrcE;
	input wire [2:0] ALUSelectE;
	input wire JumpE;
	input wire BranchSignedE;
	input wire [3:0] BSelectE;
	input wire [3:0] ZBBSelectE;
	input wire [2:0] BALUControlE;
	input wire BMUActiveE;
	input wire [1:0] CZeroE;
	output wire [1:0] FlagsE;
	output wire [$signed(P[4216-:32]) - 1:0] IEUAdrE;
	output wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcAE;
	output wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcBE;
	input wire StallM;
	input wire FlushM;
	input wire FWriteIntM;
	input wire FCvtIntW;
	input wire [$signed(P[4216-:32]) - 1:0] FIntResM;
	output wire [$signed(P[4216-:32]) - 1:0] SrcAM;
	output wire [$signed(P[4216-:32]) - 1:0] WriteDataM;
	input wire StallW;
	input wire FlushW;
	input wire RegWriteW;
	input wire IntDivW;
	input wire SquashSCW;
	input wire [2:0] ResultSrcW;
	input wire [$signed(P[4216-:32]) - 1:0] FCvtIntResW;
	input wire [$signed(P[4216-:32]) - 1:0] ReadDataW;
	input wire [$signed(P[4216-:32]) - 1:0] CSRReadValW;
	input wire [$signed(P[4216-:32]) - 1:0] MDUResultW;
	input wire [$signed(P[4216-:32]) - 1:0] FIntDivResultW;
	input wire [4:0] RdW;
	wire [$signed(P[4216-:32]) - 1:0] R1D;
	wire [$signed(P[4216-:32]) - 1:0] R2D;
	wire [$signed(P[4216-:32]) - 1:0] ImmExtD;
	wire [$signed(P[4216-:32]) - 1:0] R1E;
	wire [$signed(P[4216-:32]) - 1:0] R2E;
	wire [$signed(P[4216-:32]) - 1:0] ImmExtE;
	wire [$signed(P[4216-:32]) - 1:0] SrcAE;
	wire [$signed(P[4216-:32]) - 1:0] SrcBE;
	wire [$signed(P[4216-:32]) - 1:0] ALUResultE;
	wire [$signed(P[4216-:32]) - 1:0] AltResultE;
	wire [$signed(P[4216-:32]) - 1:0] IEUResultE;
	wire [$signed(P[4216-:32]) - 1:0] IEUResultM;
	wire [$signed(P[4216-:32]) - 1:0] IFResultM;
	wire [$signed(P[4216-:32]) - 1:0] SCResultW;
	wire [$signed(P[4216-:32]) - 1:0] ResultW;
	wire [$signed(P[4216-:32]) - 1:0] IFResultW;
	wire [$signed(P[4216-:32]) - 1:0] IFCvtResultW;
	wire [$signed(P[4216-:32]) - 1:0] MulDivResultW;
	regfile #(
		.XLEN($signed(P[4216-:32])),
		.E_SUPPORTED(P[1492])
	) regf(
		.clk(clk),
		.reset(reset),
		.we3(RegWriteW),
		.a1(Rs1D),
		.a2(Rs2D),
		.a3(RdW),
		.wd3(ResultW),
		.rd1(R1D),
		.rd2(R2D)
	);
	extend #(.P(P)) ext(
		.InstrD(InstrD[31:7]),
		.ImmSrcD(ImmSrcD),
		.ImmExtD(ImmExtD)
	);
	flopenrc #(.WIDTH($signed(P[4216-:32]))) RD1EReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(R1D),
		.q(R1E)
	);
	flopenrc #(.WIDTH($signed(P[4216-:32]))) RD2EReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(R2D),
		.q(R2E)
	);
	flopenrc #(.WIDTH($signed(P[4216-:32]))) ImmExtEReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(ImmExtD),
		.q(ImmExtE)
	);
	mux3 #(.WIDTH($signed(P[4216-:32]))) faemux(
		.d0(R1E),
		.d1(ResultW),
		.d2(IFResultM),
		.s(ForwardAE),
		.y(ForwardedSrcAE)
	);
	mux3 #(.WIDTH($signed(P[4216-:32]))) fbemux(
		.d0(R2E),
		.d1(ResultW),
		.d2(IFResultM),
		.s(ForwardBE),
		.y(ForwardedSrcBE)
	);
	comparator #(.WIDTH($signed(P[4216-:32]))) comp(
		.a(ForwardedSrcAE),
		.b(ForwardedSrcBE),
		.sgnd(BranchSignedE),
		.flags(FlagsE)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) srcamux(
		.d0(ForwardedSrcAE),
		.d1(PCE),
		.s(ALUSrcAE),
		.y(SrcAE)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) srcbmux(
		.d0(ForwardedSrcBE),
		.d1(ImmExtE),
		.s(ALUSrcBE),
		.y(SrcBE)
	);
	alu #(.P(P)) alu(
		.A(SrcAE),
		.B(SrcBE),
		.W64(W64E),
		.UW64(UW64E),
		.SubArith(SubArithE),
		.ALUSelect(ALUSelectE),
		.BSelect(BSelectE),
		.ZBBSelect(ZBBSelectE),
		.Funct3(Funct3E),
		.Funct7(Funct7E),
		.Rs2E(Rs2E),
		.BALUControl(BALUControlE),
		.BMUActive(BMUActiveE),
		.CZero(CZeroE),
		.ALUResult(ALUResultE),
		.Sum(IEUAdrE)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) altresultmux(
		.d0(ImmExtE),
		.d1(PCLinkE),
		.s(JumpE),
		.y(AltResultE)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) ieuresultmux(
		.d0(ALUResultE),
		.d1(AltResultE),
		.s(ALUResultSrcE),
		.y(IEUResultE)
	);
	flopenrc #(.WIDTH($signed(P[4216-:32]))) SrcAMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(SrcAE),
		.q(SrcAM)
	);
	flopenrc #(.WIDTH($signed(P[4216-:32]))) IEUResultMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(IEUResultE),
		.q(IEUResultM)
	);
	flopenrc #(.WIDTH($signed(P[4216-:32]))) WriteDataMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(ForwardedSrcBE),
		.q(WriteDataM)
	);
	flopenrc #(.WIDTH($signed(P[4216-:32]))) IFResultWReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(IFResultM),
		.q(IFResultW)
	);
	generate
		if (P[1491]) begin : fpmux
			mux2 #(.WIDTH($signed(P[4216-:32]))) resultmuxM(
				.d0(IEUResultM),
				.d1(FIntResM),
				.s(FWriteIntM),
				.y(IFResultM)
			);
			mux2 #(.WIDTH($signed(P[4216-:32]))) cvtresultmuxW(
				.d0(IFResultW),
				.d1(FCvtIntResW),
				.s(FCvtIntW),
				.y(IFCvtResultW)
			);
			if (P[3729] & P[1491]) begin : genblk1
				mux2 #(.WIDTH($signed(P[4216-:32]))) divresultmuxW(
					.d0(MDUResultW),
					.d1(FIntDivResultW),
					.s(IntDivW),
					.y(MulDivResultW)
				);
			end
			else begin : genblk1
				assign MulDivResultW = MDUResultW;
			end
		end
		else begin : fpmux
			assign IFResultM = IEUResultM;
			assign IFCvtResultW = IFResultW;
			assign MulDivResultW = MDUResultW;
		end
	endgenerate
	mux5 #(.WIDTH($signed(P[4216-:32]))) resultmuxW(
		.d0(IFCvtResultW),
		.d1(ReadDataW),
		.d2(CSRReadValW),
		.d3(MulDivResultW),
		.d4(SCResultW),
		.s(ResultSrcW),
		.y(ResultW)
	);
	generate
		if (P[4053]) begin : genblk2
			assign SCResultW = {{$signed(P[4216-:32]) - 1 {1'b0}}, SquashSCW};
		end
		else begin : genblk2
			assign SCResultW = 1'sb0;
		end
	endgenerate
endmodule
module extend (
	InstrD,
	ImmSrcD,
	ImmExtD
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [31:7] InstrD;
	input wire [2:0] ImmSrcD;
	output reg [$signed(P[4216-:32]) - 1:0] ImmExtD;
	localparam [$signed(P[4216-:32]) - 1:0] undefined = {$signed(P[4216-:32]) {1'bx}};
	always @(*) begin
		if (_sv2v_0)
			;
		case (ImmSrcD)
			3'b000: ImmExtD = {{$signed(P[4216-:32]) - 12 {InstrD[31]}}, InstrD[31:20]};
			3'b001: ImmExtD = {{$signed(P[4216-:32]) - 12 {InstrD[31]}}, InstrD[31:25], InstrD[11:7]};
			3'b010: ImmExtD = {{$signed(P[4216-:32]) - 12 {InstrD[31]}}, InstrD[7], InstrD[30:25], InstrD[11:8], 1'b0};
			3'b011: ImmExtD = {{$signed(P[4216-:32]) - 20 {InstrD[31]}}, InstrD[19:12], InstrD[20], InstrD[30:21], 1'b0};
			3'b100: ImmExtD = {{$signed(P[4216-:32]) - 31 {InstrD[31]}}, InstrD[30:12], 12'b000000000000};
			3'b101:
				if (((P[4053] | P[4054]) | P[4062]) | P[4061])
					ImmExtD = 1'sb0;
				else
					ImmExtD = undefined;
			default: ImmExtD = undefined;
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
module ieu (
	clk,
	reset,
	InstrD,
	STATUS_FS,
	ENVCFG_CBE,
	IllegalIEUFPUInstrD,
	IllegalBaseInstrD,
	PCE,
	PCLinkE,
	PCSrcE,
	FWriteIntE,
	FCvtIntE,
	IEUAdrE,
	IntDivE,
	W64E,
	Funct3E,
	ForwardedSrcAE,
	ForwardedSrcBE,
	RdE,
	MDUActiveE,
	CMOpM,
	IFUPrefetchE,
	LSUPrefetchM,
	SquashSCW,
	MemRWE,
	MemRWM,
	AtomicM,
	WriteDataM,
	Funct3M,
	SrcAM,
	RdM,
	FIntResM,
	InvalidateICacheM,
	FlushDCacheM,
	InstrValidD,
	InstrValidE,
	InstrValidM,
	BranchD,
	BranchE,
	JumpD,
	JumpE,
	FIntDivResultW,
	CSRReadValW,
	MDUResultW,
	FCvtIntResW,
	FCvtIntW,
	RdW,
	ReadDataW,
	StallD,
	StallE,
	StallM,
	StallW,
	FlushD,
	FlushE,
	FlushM,
	FlushW,
	StructuralStallD,
	LoadStallD,
	StoreStallD,
	CSRReadM,
	CSRWriteM,
	PrivilegedM,
	CSRWriteFenceM
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire [31:0] InstrD;
	input wire [1:0] STATUS_FS;
	input wire [3:0] ENVCFG_CBE;
	input wire IllegalIEUFPUInstrD;
	output wire IllegalBaseInstrD;
	input wire [$signed(P[4216-:32]) - 1:0] PCE;
	input wire [$signed(P[4216-:32]) - 1:0] PCLinkE;
	output wire PCSrcE;
	input wire FWriteIntE;
	input wire FCvtIntE;
	output wire [$signed(P[4216-:32]) - 1:0] IEUAdrE;
	output wire IntDivE;
	output wire W64E;
	output wire [2:0] Funct3E;
	output wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcAE;
	output wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcBE;
	output wire [4:0] RdE;
	output wire MDUActiveE;
	output wire [3:0] CMOpM;
	output wire IFUPrefetchE;
	output wire LSUPrefetchM;
	input wire SquashSCW;
	output wire [1:0] MemRWE;
	output wire [1:0] MemRWM;
	output wire [1:0] AtomicM;
	output wire [$signed(P[4216-:32]) - 1:0] WriteDataM;
	output wire [2:0] Funct3M;
	output wire [$signed(P[4216-:32]) - 1:0] SrcAM;
	output wire [4:0] RdM;
	input wire [$signed(P[4216-:32]) - 1:0] FIntResM;
	output wire InvalidateICacheM;
	output wire FlushDCacheM;
	output wire InstrValidD;
	output wire InstrValidE;
	output wire InstrValidM;
	output wire BranchD;
	output wire BranchE;
	output wire JumpD;
	output wire JumpE;
	input wire [$signed(P[4216-:32]) - 1:0] FIntDivResultW;
	input wire [$signed(P[4216-:32]) - 1:0] CSRReadValW;
	input wire [$signed(P[4216-:32]) - 1:0] MDUResultW;
	input wire [$signed(P[4216-:32]) - 1:0] FCvtIntResW;
	input wire FCvtIntW;
	output wire [4:0] RdW;
	input wire [$signed(P[4216-:32]) - 1:0] ReadDataW;
	input wire StallD;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushD;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	output wire StructuralStallD;
	output wire LoadStallD;
	output wire StoreStallD;
	output wire CSRReadM;
	output wire CSRWriteM;
	output wire PrivilegedM;
	output wire CSRWriteFenceM;
	wire [2:0] ImmSrcD;
	wire [1:0] FlagsE;
	wire ALUSrcAE;
	wire ALUSrcBE;
	wire [2:0] ResultSrcW;
	wire ALUResultSrcE;
	wire [2:0] ALUSelectE;
	wire FWriteIntM;
	wire IntDivW;
	wire [3:0] BSelectE;
	wire [3:0] ZBBSelectE;
	wire [2:0] BALUControlE;
	wire SubArithE;
	wire UW64E;
	wire [6:0] Funct7E;
	wire [4:0] Rs1D;
	wire [4:0] Rs2D;
	wire [4:0] Rs2E;
	wire [1:0] ForwardAE;
	wire [1:0] ForwardBE;
	wire RegWriteW;
	wire BranchSignedE;
	wire BMUActiveE;
	wire [1:0] CZeroE;
	controller #(.P(P)) c(
		.clk(clk),
		.reset(reset),
		.StallD(StallD),
		.FlushD(FlushD),
		.InstrD(InstrD),
		.STATUS_FS(STATUS_FS),
		.ENVCFG_CBE(ENVCFG_CBE),
		.ImmSrcD(ImmSrcD),
		.IllegalIEUFPUInstrD(IllegalIEUFPUInstrD),
		.IllegalBaseInstrD(IllegalBaseInstrD),
		.StructuralStallD(StructuralStallD),
		.LoadStallD(LoadStallD),
		.StoreStallD(StoreStallD),
		.Rs1D(Rs1D),
		.Rs2D(Rs2D),
		.Rs2E(Rs2E),
		.StallE(StallE),
		.FlushE(FlushE),
		.FlagsE(FlagsE),
		.FWriteIntE(FWriteIntE),
		.PCSrcE(PCSrcE),
		.ALUSrcAE(ALUSrcAE),
		.ALUSrcBE(ALUSrcBE),
		.ALUResultSrcE(ALUResultSrcE),
		.ALUSelectE(ALUSelectE),
		.Funct3E(Funct3E),
		.Funct7E(Funct7E),
		.IntDivE(IntDivE),
		.W64E(W64E),
		.UW64E(UW64E),
		.SubArithE(SubArithE),
		.BranchD(BranchD),
		.BranchE(BranchE),
		.JumpD(JumpD),
		.JumpE(JumpE),
		.BranchSignedE(BranchSignedE),
		.BSelectE(BSelectE),
		.ZBBSelectE(ZBBSelectE),
		.BALUControlE(BALUControlE),
		.BMUActiveE(BMUActiveE),
		.CZeroE(CZeroE),
		.MDUActiveE(MDUActiveE),
		.FCvtIntE(FCvtIntE),
		.ForwardAE(ForwardAE),
		.ForwardBE(ForwardBE),
		.CMOpM(CMOpM),
		.IFUPrefetchE(IFUPrefetchE),
		.LSUPrefetchM(LSUPrefetchM),
		.StallM(StallM),
		.FlushM(FlushM),
		.MemRWE(MemRWE),
		.MemRWM(MemRWM),
		.CSRReadM(CSRReadM),
		.CSRWriteM(CSRWriteM),
		.PrivilegedM(PrivilegedM),
		.AtomicM(AtomicM),
		.Funct3M(Funct3M),
		.FlushDCacheM(FlushDCacheM),
		.InstrValidM(InstrValidM),
		.InstrValidE(InstrValidE),
		.InstrValidD(InstrValidD),
		.FWriteIntM(FWriteIntM),
		.StallW(StallW),
		.FlushW(FlushW),
		.RegWriteW(RegWriteW),
		.IntDivW(IntDivW),
		.ResultSrcW(ResultSrcW),
		.CSRWriteFenceM(CSRWriteFenceM),
		.InvalidateICacheM(InvalidateICacheM),
		.RdW(RdW),
		.RdE(RdE),
		.RdM(RdM)
	);
	datapath #(.P(P)) dp(
		.clk(clk),
		.reset(reset),
		.ImmSrcD(ImmSrcD),
		.InstrD(InstrD),
		.Rs1D(Rs1D),
		.Rs2D(Rs2D),
		.Rs2E(Rs2E),
		.StallE(StallE),
		.FlushE(FlushE),
		.ForwardAE(ForwardAE),
		.ForwardBE(ForwardBE),
		.W64E(W64E),
		.UW64E(UW64E),
		.SubArithE(SubArithE),
		.Funct3E(Funct3E),
		.Funct7E(Funct7E),
		.ALUSrcAE(ALUSrcAE),
		.ALUSrcBE(ALUSrcBE),
		.ALUResultSrcE(ALUResultSrcE),
		.ALUSelectE(ALUSelectE),
		.JumpE(JumpE),
		.BranchSignedE(BranchSignedE),
		.PCE(PCE),
		.PCLinkE(PCLinkE),
		.FlagsE(FlagsE),
		.IEUAdrE(IEUAdrE),
		.ForwardedSrcAE(ForwardedSrcAE),
		.ForwardedSrcBE(ForwardedSrcBE),
		.BSelectE(BSelectE),
		.ZBBSelectE(ZBBSelectE),
		.BALUControlE(BALUControlE),
		.BMUActiveE(BMUActiveE),
		.CZeroE(CZeroE),
		.StallM(StallM),
		.FlushM(FlushM),
		.FWriteIntM(FWriteIntM),
		.FIntResM(FIntResM),
		.SrcAM(SrcAM),
		.WriteDataM(WriteDataM),
		.FCvtIntW(FCvtIntW),
		.StallW(StallW),
		.FlushW(FlushW),
		.RegWriteW(RegWriteW),
		.IntDivW(IntDivW),
		.SquashSCW(SquashSCW),
		.ResultSrcW(ResultSrcW),
		.ReadDataW(ReadDataW),
		.FCvtIntResW(FCvtIntResW),
		.CSRReadValW(CSRReadValW),
		.MDUResultW(MDUResultW),
		.FIntDivResultW(FIntDivResultW),
		.RdW(RdW)
	);
endmodule
module regfile (
	clk,
	reset,
	we3,
	a1,
	a2,
	a3,
	wd3,
	rd1,
	rd2
);
	parameter XLEN = 0;
	parameter E_SUPPORTED = 0;
	input wire clk;
	input wire reset;
	input wire we3;
	input wire [4:0] a1;
	input wire [4:0] a2;
	input wire [4:0] a3;
	input wire [XLEN - 1:0] wd3;
	output wire [XLEN - 1:0] rd1;
	output wire [XLEN - 1:0] rd2;
	localparam NUMREGS = (E_SUPPORTED ? 16 : 32);
	reg [XLEN - 1:0] rf [NUMREGS - 1:1];
	integer i;
	always @(negedge clk)
		if (reset)
			for (i = 1; i < NUMREGS; i = i + 1)
				rf[i] <= 1'sb0;
		else if (we3)
			rf[a3] <= wd3;
	assign rd1 = (a1 != 0 ? rf[a1] : 0);
	assign rd2 = (a2 != 0 ? rf[a2] : 0);
endmodule
module shifter (
	A,
	Amt,
	Right,
	Rotate,
	W64,
	SubArith,
	Y
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[4216-:32]) - 1:0] A;
	input wire [$signed(P[1485-:32]) - 1:0] Amt;
	input wire Right;
	input wire Rotate;
	input wire W64;
	input wire SubArith;
	output wire [$signed(P[4216-:32]) - 1:0] Y;
	reg [(2 * $signed(P[4216-:32])) - 2:0] Z;
	wire [(2 * $signed(P[4216-:32])) - 2:0] ZShift;
	wire [$signed(P[1485-:32]) - 1:0] TruncAmt;
	wire [$signed(P[1485-:32]) - 1:0] Offset;
	wire Sign;
	assign Sign = A[$signed(P[4216-:32]) - 1] & SubArith;
	generate
		if ($signed(P[4216-:32]) == 32) begin : genblk1
			if (P[1757] | P[1750]) begin : rotfunnel32
				always @(*) begin
					if (_sv2v_0)
						;
					case ({Right, Rotate})
						2'b00: Z = {A[31:0], 31'b0000000000000000000000000000000};
						2'b01: Z = {A[31:0], A[31:1]};
						2'b10: Z = {{31 {Sign}}, A[31:0]};
						2'b11: Z = {A[30:0], A[31:0]};
					endcase
				end
			end
			else begin : norotfunnel32
				always @(*) begin
					if (_sv2v_0)
						;
					if (Right)
						Z = {{31 {Sign}}, A[31:0]};
					else
						Z = {A[31:0], 31'b0000000000000000000000000000000};
				end
			end
			assign TruncAmt = Amt;
		end
		else begin : genblk1
			wire [$signed(P[4216-:32]) - 1:0] A64;
			mux3 #(.WIDTH(64)) extendmux(
				.d0({{32 {1'b0}}, A[31:0]}),
				.d1({{32 {A[31]}}, A[31:0]}),
				.d2(A),
				.s({~W64, SubArith}),
				.y(A64)
			);
			if (P[1757] | P[1750]) begin : rotfunnel64
				wire [$signed(P[4216-:32]) - 1:0] RotA;
				mux2 #(.WIDTH($signed(P[4216-:32]))) rotmux(
					.d0(A),
					.d1({A[31:0], A[31:0]}),
					.s(W64),
					.y(RotA)
				);
				always @(*) begin
					if (_sv2v_0)
						;
					case ({Right, Rotate})
						2'b00: Z = {A64[63:0], 63'b000000000000000000000000000000000000000000000000000000000000000};
						2'b01: Z = {RotA[63:0], RotA[63:1]};
						2'b10: Z = {{63 {Sign}}, A64[63:0]};
						2'b11: Z = {RotA[62:0], RotA[63:0]};
					endcase
				end
			end
			else begin : norotfunnel64
				always @(*) begin
					if (_sv2v_0)
						;
					if (Right)
						Z = {{63 {Sign}}, A64[63:0]};
					else
						Z = {A64[63:0], 63'b000000000000000000000000000000000000000000000000000000000000000};
				end
			end
			assign TruncAmt = (W64 ? {1'b0, Amt[4:0]} : Amt);
		end
	endgenerate
	assign Offset = (Right ? TruncAmt : ~TruncAmt);
	assign ZShift = Z >> Offset;
	assign Y = ZShift[$signed(P[4216-:32]) - 1:0];
	initial _sv2v_0 = 0;
endmodule
module decompress (
	InstrRawD,
	InstrD,
	IllegalCompInstrD
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [31:0] InstrRawD;
	output wire [31:0] InstrD;
	output wire IllegalCompInstrD;
	reg [32:0] LInstrD;
	wire [15:0] instr16;
	wire [4:0] rds1;
	wire [4:0] rs2;
	wire [4:0] rs1p;
	wire [4:0] rs2p;
	wire [4:0] rds1p;
	wire [4:0] rdp;
	wire [11:0] immCILSP;
	wire [11:0] immCILSPD;
	wire [11:0] immCSS;
	wire [11:0] immCSSD;
	wire [11:0] immCL;
	wire [11:0] immCLD;
	wire [11:0] immCI;
	wire [11:0] immCS;
	wire [11:0] immCSD;
	wire [11:0] immCB;
	wire [11:0] immCIASP;
	wire [11:0] immCIW;
	wire [19:0] immCJ;
	wire [19:0] immCILUI;
	wire [5:0] immSH;
	wire [1:0] op;
	wire LegalCompInstrD;
	assign instr16 = InstrRawD[15:0];
	assign op = instr16[1:0];
	assign rds1 = instr16[11:7];
	assign rs2 = instr16[6:2];
	assign rs1p = {2'b01, instr16[9:7]};
	assign rds1p = {2'b01, instr16[9:7]};
	assign rs2p = {2'b01, instr16[4:2]};
	assign rdp = {2'b01, instr16[4:2]};
	assign immCILSP = {4'b0000, instr16[3:2], instr16[12], instr16[6:4], 2'b00};
	assign immCILSPD = {3'b000, instr16[4:2], instr16[12], instr16[6:5], 3'b000};
	assign immCSS = {4'b0000, instr16[8:7], instr16[12:9], 2'b00};
	assign immCSSD = {3'b000, instr16[9:7], instr16[12:10], 3'b000};
	assign immCL = {5'b00000, instr16[5], instr16[12:10], instr16[6], 2'b00};
	assign immCLD = {4'b0000, instr16[6:5], instr16[12:10], 3'b000};
	assign immCS = {5'b00000, instr16[5], instr16[12:10], instr16[6], 2'b00};
	assign immCSD = {4'b0000, instr16[6:5], instr16[12:10], 3'b000};
	assign immCJ = {instr16[12], instr16[8], instr16[10:9], instr16[6], instr16[7], instr16[2], instr16[11], instr16[5:3], {9 {instr16[12]}}};
	assign immCB = {{4 {instr16[12]}}, instr16[6:5], instr16[2], instr16[11:10], instr16[4:3], instr16[12]};
	assign immCI = {{7 {instr16[12]}}, instr16[6:2]};
	assign immCILUI = {{15 {instr16[12]}}, instr16[6:2]};
	assign immCIASP = {{3 {instr16[12]}}, instr16[4:3], instr16[5], instr16[2], instr16[6], 4'b0000};
	assign immCIW = {2'b00, instr16[10:7], instr16[12:11], instr16[5], instr16[6], 2'b00};
	assign immSH = {instr16[12], instr16[6:2]};
	always @(*) begin
		if (_sv2v_0)
			;
		if (op == 2'b11)
			LInstrD = {1'b1, InstrRawD};
		else begin
			LInstrD = {17'b00000000000000000, instr16};
			case ({op, instr16[15:13]})
				5'b00000:
					if (immCIW != 0)
						LInstrD = {1'b1, immCIW, 8'b00010000, rdp, 7'b0010011};
				5'b00001:
					if (P[1752])
						LInstrD = {1'b1, immCLD, rs1p, 3'b011, rdp, 7'b0000111};
				5'b00010: LInstrD = {1'b1, immCL, rs1p, 3'b010, rdp, 7'b0000011};
				5'b00011:
					if ($signed(P[4216-:32]) == 32) begin
						if (P[1751])
							LInstrD = {1'b1, immCL, rs1p, 3'b010, rdp, 7'b0000111};
					end
					else
						LInstrD = {1'b1, immCLD, rs1p, 3'b011, rdp, 7'b0000011};
				5'b00100:
					if (P[1753]) begin
						if (instr16[12:10] == 3'b000)
							LInstrD = {11'b10000000000, instr16[5], instr16[6], rs1p, 3'b100, rdp, 7'b0000011};
						else if (instr16[12:10] == 3'b001) begin
							if (instr16[6])
								LInstrD = {11'b10000000000, instr16[5], 1'b0, rs1p, 3'b001, rdp, 7'b0000011};
							else
								LInstrD = {11'b10000000000, instr16[5], 1'b0, rs1p, 3'b101, rdp, 7'b0000011};
						end
						else if (instr16[12:10] == 3'b010)
							LInstrD = {8'b10000000, rs2p, rs1p, 6'b000000, instr16[5], instr16[6], 7'b0100011};
						else if ((instr16[12:10] == 3'b011) & (instr16[6] == 1'b0))
							LInstrD = {8'b10000000, rs2p, rs1p, 6'b001000, instr16[5], 8'b00100011};
					end
				5'b00101:
					if (P[1752])
						LInstrD = {1'b1, immCSD[11:5], rs2p, rs1p, 3'b011, immCSD[4:0], 7'b0100111};
				5'b00110: LInstrD = {1'b1, immCS[11:5], rs2p, rs1p, 3'b010, immCS[4:0], 7'b0100011};
				5'b00111:
					if ($signed(P[4216-:32]) == 32) begin
						if (P[1751])
							LInstrD = {1'b1, immCS[11:5], rs2p, rs1p, 3'b010, immCS[4:0], 7'b0100111};
					end
					else
						LInstrD = {1'b1, immCSD[11:5], rs2p, rs1p, 3'b011, immCSD[4:0], 7'b0100011};
				5'b01000:
					if (rds1 != 5'b00000) begin
						if (immCI[5:0] != 0)
							LInstrD = {1'b1, immCI, rds1, 3'b000, rds1, 7'b0010011};
						else
							LInstrD = 33'b100000000000000000000000000010011;
					end
					else if (immCI[5:0] == 6'b000000)
						LInstrD = 33'b100000000000000000000000000010011;
					else
						LInstrD = 33'b100000000000000000000000000010011;
				5'b01001:
					if ($signed(P[4216-:32]) == 32)
						LInstrD = {1'b1, immCJ, 12'b000011101111};
					else if (rds1 != 5'b00000)
						LInstrD = {1'b1, immCI, rds1, 3'b000, rds1, 7'b0011011};
				5'b01010:
					if (rds1 != 5'b00000)
						LInstrD = {1'b1, immCI, 8'b00000000, rds1, 7'b0010011};
					else
						LInstrD = 33'b100000000000000000000000000010011;
				5'b01011:
					if (rds1 == 5'b00010) begin
						if (immCIASP[9:4] != 6'b000000)
							LInstrD = {1'b1, immCIASP, rds1, 3'b000, rds1, 7'b0010011};
					end
					else if (immCILUI[5:0] != 0) begin
						if (rds1 != 5'b00000)
							LInstrD = {1'b1, immCILUI, rds1, 7'b0110111};
						else
							LInstrD = 33'b100000000000000000000000000010011;
					end
				5'b01100:
					if (instr16[11:10] == 2'b00) begin
						if (($signed(P[4216-:32]) > 32) | ~immSH[5])
							LInstrD = {7'b1000000, immSH, rds1p, 3'b101, rds1p, 7'b0010011};
					end
					else if (instr16[11:10] == 2'b01) begin
						if (($signed(P[4216-:32]) > 32) | ~immSH[5])
							LInstrD = {7'b1010000, immSH, rds1p, 3'b101, rds1p, 7'b0010011};
					end
					else if (instr16[11:10] == 2'b10)
						LInstrD = {1'b1, immCI, rds1p, 3'b111, rds1p, 7'b0010011};
					else if (instr16[12:10] == 3'b011) begin
						if (instr16[6:5] == 2'b00)
							LInstrD = {8'b10100000, rs2p, rds1p, 3'b000, rds1p, 7'b0110011};
						else if (instr16[6:5] == 2'b01)
							LInstrD = {8'b10000000, rs2p, rds1p, 3'b100, rds1p, 7'b0110011};
						else if (instr16[6:5] == 2'b10)
							LInstrD = {8'b10000000, rs2p, rds1p, 3'b110, rds1p, 7'b0110011};
						else
							LInstrD = {8'b10000000, rs2p, rds1p, 3'b111, rds1p, 7'b0110011};
					end
					else if ((instr16[6:5] == 2'b00) & ($signed(P[4216-:32]) > 32))
						LInstrD = {8'b10100000, rs2p, rds1p, 3'b000, rds1p, 7'b0111011};
					else if ((instr16[6:5] == 2'b01) & ($signed(P[4216-:32]) > 32))
						LInstrD = {8'b10000000, rs2p, rds1p, 3'b000, rds1p, 7'b0111011};
					else if ((instr16[6:2] == 5'b11000) & P[1753])
						LInstrD = {13'b1000011111111, rds1p, 3'b111, rds1p, 7'b0010011};
					else if (((instr16[6:2] == 5'b11001) & P[1753]) & P[1757])
						LInstrD = {13'b1011000000100, rds1p, 3'b001, rds1p, 7'b0010011};
					else if (((instr16[6:2] == 5'b11010) & P[1753]) & P[1757])
						LInstrD = {13'b1000010000000, rds1p, 3'b100, rds1p, 3'b011, $signed(P[4216-:32]) > 32, 3'b011};
					else if (((instr16[6:2] == 5'b11011) & P[1753]) & P[1757])
						LInstrD = {13'b1011000000101, rds1p, 3'b001, rds1p, 7'b0010011};
					else if ((instr16[6:2] == 5'b11101) & P[1753])
						LInstrD = {13'b1111111111111, rds1p, 3'b100, rds1p, 7'b0010011};
					else if ((((instr16[6:2] == 5'b11100) & P[1753]) & P[1758]) & ($signed(P[4216-:32]) > 32))
						LInstrD = {13'b1000010000000, rds1p, 3'b000, rds1p, 7'b0111011};
					else if (((instr16[6:5] == 2'b10) & P[1753]) & P[4063])
						LInstrD = {8'b10000001, rs2p, rds1p, 3'b000, rds1p, 7'b0110011};
				5'b01101: LInstrD = {1'b1, immCJ, 12'b000001101111};
				5'b01110: LInstrD = {1'b1, immCB[11:5], 5'b00000, rs1p, 3'b000, immCB[4:0], 7'b1100011};
				5'b01111: LInstrD = {1'b1, immCB[11:5], 5'b00000, rs1p, 3'b001, immCB[4:0], 7'b1100011};
				5'b10000:
					if (immSH != 0) begin
						if (($signed(P[4216-:32]) > 32) | ~immSH[5]) begin
							if (rds1 != 5'b00000)
								LInstrD = {7'b1000000, immSH, rds1, 3'b001, rds1, 7'b0010011};
							else
								LInstrD = 33'b100000000000000000000000000010011;
						end
					end
					else
						LInstrD = 33'b100000000000000000000000000010011;
				5'b10001:
					if (P[1752])
						LInstrD = {1'b1, immCILSPD, 8'b00010011, rds1, 7'b0000111};
				5'b10010:
					if (rds1 != 5'b00000)
						LInstrD = {1'b1, immCILSP, 8'b00010010, rds1, 7'b0000011};
				5'b10011:
					if ($signed(P[4216-:32]) == 32) begin
						if (P[1751])
							LInstrD = {1'b1, immCILSP, 8'b00010010, rds1, 7'b0000111};
					end
					else if (rds1 != 5'b00000)
						LInstrD = {1'b1, immCILSPD, 8'b00010011, rds1, 7'b0000011};
				5'b10100:
					if (instr16[12] == 0) begin
						if (rs2 == 5'b00000) begin
							if (rds1 != 5'b00000)
								LInstrD = {13'b1000000000000, rds1, 15'b000000001100111};
						end
						else if (rds1 != 5'b00000)
							LInstrD = {8'b10000000, rs2, 8'b00000000, rds1, 7'b0110011};
						else
							LInstrD = 33'b100000000000000000000000000010011;
					end
					else if (rs2 == 5'b00000) begin
						if (rds1 == 5'b00000)
							LInstrD = 33'b100000000000100000000000001110011;
						else
							LInstrD = {13'b1000000000000, rds1, 15'b000000011100111};
					end
					else if (rds1 != 0)
						LInstrD = {8'b10000000, rs2, rds1, 3'b000, rds1, 7'b0110011};
					else
						LInstrD = 33'b100000000000000000000000000010011;
				5'b10101:
					if (P[1752])
						LInstrD = {1'b1, immCSSD[11:5], rs2, 8'b00010011, immCSSD[4:0], 7'b0100111};
				5'b10110: LInstrD = {1'b1, immCSS[11:5], rs2, 8'b00010010, immCSS[4:0], 7'b0100011};
				5'b10111:
					if ($signed(P[4216-:32]) == 32) begin
						if (P[1751])
							LInstrD = {1'b1, immCSS[11:5], rs2, 8'b00010010, immCSS[4:0], 7'b0100111};
					end
					else
						LInstrD = {1'b1, immCSSD[11:5], rs2, 8'b00010011, immCSSD[4:0], 7'b0100011};
				default:
					;
			endcase
		end
	end
	assign {LegalCompInstrD, InstrD} = LInstrD;
	assign IllegalCompInstrD = ~LegalCompInstrD;
	initial _sv2v_0 = 0;
endmodule
module ifu (
	clk,
	reset,
	StallF,
	StallD,
	StallE,
	StallM,
	StallW,
	FlushD,
	FlushE,
	FlushM,
	FlushW,
	IFUStallF,
	InvalidateICacheM,
	CSRWriteFenceM,
	InstrValidD,
	InstrValidE,
	BranchD,
	BranchE,
	JumpD,
	JumpE,
	IFUHADDR,
	HRDATA,
	IFUHREADY,
	IFUHWRITE,
	IFUHSIZE,
	IFUHBURST,
	IFUHTRANS,
	PCSpillF,
	PCLinkE,
	PCSrcE,
	IEUAdrE,
	IEUAdrM,
	PCE,
	BPWrongE,
	BPWrongM,
	CommittedF,
	EPCM,
	TrapVectorM,
	RetM,
	TrapM,
	InstrD,
	InstrM,
	InstrOrigM,
	PCM,
	IClassM,
	BPDirWrongM,
	BTAWrongM,
	RASPredPCWrongM,
	IClassWrongM,
	ICacheStallF,
	IllegalBaseInstrD,
	IllegalFPUInstrD,
	InstrPageFaultF,
	IllegalIEUFPUInstrD,
	InstrMisalignedFaultM,
	PrivilegeModeW,
	PTE,
	PageType,
	ITLBWriteF,
	SATP_REGW,
	STATUS_MXR,
	STATUS_SUM,
	STATUS_MPRV,
	STATUS_MPP,
	ENVCFG_PBMTE,
	ENVCFG_ADUE,
	sfencevmaM,
	ITLBMissOrUpdateAF,
	PMPCFG_ARRAY_REGW,
	PMPADDR_ARRAY_REGW,
	InstrAccessFaultF,
	ICacheAccess,
	ICacheMiss
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallF;
	input wire StallD;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushD;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	output wire IFUStallF;
	input wire InvalidateICacheM;
	input wire CSRWriteFenceM;
	input wire InstrValidD;
	input wire InstrValidE;
	input wire BranchD;
	input wire BranchE;
	input wire JumpD;
	input wire JumpE;
	output wire [$signed(P[1640-:32]) - 1:0] IFUHADDR;
	input wire [$signed(P[4216-:32]) - 1:0] HRDATA;
	input wire IFUHREADY;
	output wire IFUHWRITE;
	output wire [2:0] IFUHSIZE;
	output wire [2:0] IFUHBURST;
	output wire [1:0] IFUHTRANS;
	output wire [$signed(P[4216-:32]) - 1:0] PCSpillF;
	output wire [$signed(P[4216-:32]) - 1:0] PCLinkE;
	input wire PCSrcE;
	input wire [$signed(P[4216-:32]) - 1:0] IEUAdrE;
	input wire [$signed(P[4216-:32]) - 1:0] IEUAdrM;
	output wire [$signed(P[4216-:32]) - 1:0] PCE;
	output wire BPWrongE;
	output wire BPWrongM;
	output wire CommittedF;
	input wire [$signed(P[4216-:32]) - 1:0] EPCM;
	input wire [$signed(P[4216-:32]) - 1:0] TrapVectorM;
	input wire RetM;
	input wire TrapM;
	output wire [31:0] InstrD;
	output wire [31:0] InstrM;
	output wire [31:0] InstrOrigM;
	output wire [$signed(P[4216-:32]) - 1:0] PCM;
	output wire [3:0] IClassM;
	output wire BPDirWrongM;
	output wire BTAWrongM;
	output wire RASPredPCWrongM;
	output wire IClassWrongM;
	output wire ICacheStallF;
	input wire IllegalBaseInstrD;
	input wire IllegalFPUInstrD;
	output wire InstrPageFaultF;
	output wire IllegalIEUFPUInstrD;
	output wire InstrMisalignedFaultM;
	input wire [1:0] PrivilegeModeW;
	input wire [$signed(P[4216-:32]) - 1:0] PTE;
	input wire [1:0] PageType;
	input wire ITLBWriteF;
	input wire [$signed(P[4216-:32]) - 1:0] SATP_REGW;
	input wire STATUS_MXR;
	input wire STATUS_SUM;
	input wire STATUS_MPRV;
	input wire [1:0] STATUS_MPP;
	input wire ENVCFG_PBMTE;
	input wire ENVCFG_ADUE;
	input wire sfencevmaM;
	output wire ITLBMissOrUpdateAF;
	input wire [($signed(P[3728-:32]) * 8) - 1:0] PMPCFG_ARRAY_REGW;
	input wire [(($signed(P[1640-:32]) - 3) >= 0 ? ($signed(P[3728-:32]) * ($signed(P[1640-:32]) - 2)) - 1 : ($signed(P[3728-:32]) * (4 - $signed(P[1640-:32]))) + ($signed(P[1640-:32]) - 4)):(($signed(P[1640-:32]) - 3) >= 0 ? 0 : $signed(P[1640-:32]) - 3)] PMPADDR_ARRAY_REGW;
	output wire InstrAccessFaultF;
	output wire ICacheAccess;
	output wire ICacheMiss;
	localparam [31:0] nop = 32'h00000013;
	localparam LINELEN = (P[4050] ? $signed(P[3825-:32]) : $signed(P[4216-:32]));
	wire [$signed(P[4216-:32]) - 1:0] PCNextF;
	wire [$signed(P[4216-:32]) - 1:0] PC1NextF;
	wire [$signed(P[4216-:32]) - 1:0] PC2NextF;
	wire [$signed(P[4216-:32]) - 1:0] UnalignedPCNextF;
	wire BranchMisalignedFaultE;
	reg [$signed(P[4216-:32]) - 1:0] PCPlus2or4F;
	wire [$signed(P[4216-:32]) - 1:0] PCSpillNextF;
	wire [$signed(P[4216-:32]) - 1:2] PCPlus4F;
	wire [$signed(P[4216-:32]) - 1:0] PCD;
	wire [$signed(P[4216-:32]) - 1:0] NextValidPCE;
	wire [$signed(P[4216-:32]) - 1:0] PCF;
	wire [$signed(P[1640-:32]) - 1:0] PCPF;
	wire [$signed(P[4216-:32]) + 1:0] PCFExt;
	wire [31:0] IROMInstrF;
	wire [31:0] ICacheInstrF;
	wire [31:0] InstrRawF;
	wire CompressedF;
	wire CompressedE;
	wire [31:0] PostSpillInstrRawF;
	wire [31:0] InstrRawD;
	wire IllegalIEUInstrD;
	wire [1:0] IFURWF;
	wire [31:0] InstrE;
	wire [31:0] NextInstrD;
	wire [31:0] NextInstrE;
	wire CacheableF;
	wire SelSpillNextF;
	wire BusStall;
	wire IFUCacheBusStallF;
	wire GatedStallD;
	wire BusCommittedF;
	wire CacheCommittedF;
	wire SelIROM;
	wire [15:0] InstrRawE;
	wire [15:0] InstrRawM;
	wire [LINELEN - 1:0] FetchBuffer;
	wire [31:0] ShiftUncachedInstr;
	wire ITLBMissF;
	wire InstrUpdateAF;
	assign PCFExt = {2'b00, PCSpillF};
	generate
		if (P[1754]) begin : Spill
			spill #(.P(P)) spill(
				.clk(clk),
				.reset(reset),
				.StallF(StallF),
				.FlushD(FlushD),
				.PCF(PCF),
				.PCPlus4F(PCPlus4F),
				.PCNextF(PCNextF),
				.InstrRawF(InstrRawF),
				.CacheableF(CacheableF),
				.IFUCacheBusStallF(IFUCacheBusStallF),
				.ITLBMissOrUpdateAF(ITLBMissOrUpdateAF),
				.PCSpillNextF(PCSpillNextF),
				.PCSpillF(PCSpillF),
				.SelSpillNextF(SelSpillNextF),
				.PostSpillInstrRawF(PostSpillInstrRawF),
				.CompressedF(CompressedF)
			);
		end
		else begin : NoSpill
			assign PCSpillNextF = PCNextF;
			assign PCSpillF = PCF;
			assign PostSpillInstrRawF = InstrRawF;
			assign {SelSpillNextF, CompressedF} = 1'sb0;
		end
		if (P[4086] == 1) begin : immu
			wire StallMQ;
			wire TLBFlush;
			flopr #(.WIDTH(1)) StallMReg(
				.clk(clk),
				.reset(reset),
				.d(StallM),
				.q(StallMQ)
			);
			assign TLBFlush = sfencevmaM & ~StallMQ;
			mmu #(
				.P(P),
				.TLB_ENTRIES($signed(P[4049-:32])),
				.IMMU(1)
			) immu(
				.clk(clk),
				.reset(reset),
				.SATP_REGW(SATP_REGW),
				.STATUS_MXR(STATUS_MXR),
				.STATUS_SUM(STATUS_SUM),
				.STATUS_MPRV(STATUS_MPRV),
				.STATUS_MPP(STATUS_MPP),
				.ENVCFG_PBMTE(ENVCFG_PBMTE),
				.ENVCFG_ADUE(ENVCFG_ADUE),
				.PrivilegeModeW(PrivilegeModeW),
				.DisableTranslation(1'b0),
				.VAdr(PCFExt),
				.Size(2'b10),
				.PTE(PTE),
				.PageTypeWriteVal(PageType),
				.TLBWrite(ITLBWriteF),
				.TLBFlush(TLBFlush),
				.PhysicalAddress(PCPF),
				.TLBMiss(ITLBMissF),
				.Cacheable(CacheableF),
				.Idempotent(),
				.SelTIM(SelIROM),
				.InstrAccessFaultF(InstrAccessFaultF),
				.LoadAccessFaultM(),
				.StoreAmoAccessFaultM(),
				.InstrPageFaultF(InstrPageFaultF),
				.LoadPageFaultM(),
				.StoreAmoPageFaultM(),
				.LoadMisalignedFaultM(),
				.StoreAmoMisalignedFaultM(),
				.UpdateDA(InstrUpdateAF),
				.CMOpM(4'b0000),
				.AtomicAccessM(1'b0),
				.ExecuteAccessF(1'b1),
				.WriteAccessM(1'b0),
				.ReadAccessM(1'b0),
				.PMPCFG_ARRAY_REGW(PMPCFG_ARRAY_REGW),
				.PMPADDR_ARRAY_REGW(PMPADDR_ARRAY_REGW)
			);
			assign ITLBMissOrUpdateAF = ITLBMissF | (P[4064] & InstrUpdateAF);
		end
		else begin : genblk2
			assign {ITLBMissF, InstrAccessFaultF, InstrPageFaultF, InstrUpdateAF} = 1'sb0;
			assign PCPF = PCFExt[$signed(P[1640-:32]) - 1:0];
			assign CacheableF = 1'b1;
			assign SelIROM = 1'sb0;
			assign ITLBMissOrUpdateAF = 1'sb0;
		end
	endgenerate
	assign CommittedF = CacheCommittedF | BusCommittedF;
	generate
		if (P[3471]) begin : irom
			wire IROMce;
			assign IROMce = ~GatedStallD | reset;
			assign IFURWF = 2'b10;
			irom #(.P(P)) irom(
				.clk(clk),
				.ce(IROMce),
				.Adr(PCSpillNextF[$signed(P[4216-:32]) - 1:0]),
				.IROMInstrF(IROMInstrF)
			);
		end
		else begin : genblk3
			assign IFURWF = 2'b10;
			assign IROMInstrF = 1'sb0;
		end
		if (P[4052]) begin : bus
			localparam BEATSPERLINE = (P[4050] ? $signed(P[3825-:32]) / $signed(P[4151-:32]) : 1);
			localparam AHBWLOGBWPL = (P[4050] ? $clog2(BEATSPERLINE) : 1);
			if (P[4050]) begin : icache
				localparam LLENPOVERAHBW = $signed(P[383-:32]) / $signed(P[4151-:32]);
				wire [$signed(P[1640-:32]) - 1:0] ICacheBusAdr;
				wire ICacheBusAck;
				wire [1:0] CacheBusRW;
				wire [1:0] BusRW;
				wire [1:0] CacheRWF;
				assign BusRW = ((~ITLBMissF & ~CacheableF) & ~SelIROM ? IFURWF : {2 {1'sb0}});
				assign CacheRWF = ((~ITLBMissF & CacheableF) & ~SelIROM ? IFURWF : {2 {1'sb0}});
				localparam [0:0] sv2v_uu_icache_ext_SelHPTW_0 = 1'sb0;
				localparam sv2v_uu_icache_WORDLEN = 32;
				localparam [3:0] sv2v_uu_icache_ext_ByteMask_0 = 1'sb0;
				localparam sv2v_uu_icache_LOGBWPL = AHBWLOGBWPL;
				localparam [sv2v_uu_icache_LOGBWPL - 1:0] sv2v_uu_icache_ext_BeatCount_0 = 1'sb0;
				localparam [0:0] sv2v_uu_icache_ext_SelBusBeat_0 = 1'sb0;
				localparam [31:0] sv2v_uu_icache_ext_WriteData_0 = 1'sb0;
				localparam [0:0] sv2v_uu_icache_ext_FlushCache_0 = 1'sb0;
				localparam [3:0] sv2v_uu_icache_ext_CMOpM_0 = 1'sb0;
				cache #(
					.P(P),
					.PA_BITS($signed(P[1640-:32])),
					.LINELEN($signed(P[3825-:32])),
					.NUMSETS(($signed(P[3857-:32]) * 8) / $signed(P[3825-:32])),
					.NUMWAYS($signed(P[3889-:32])),
					.LOGBWPL(AHBWLOGBWPL),
					.WORDLEN(32),
					.MUXINTERVAL(16),
					.READ_ONLY_CACHE(1)
				) icache(
					.clk(clk),
					.reset(reset),
					.FlushStage(FlushD),
					.Stall(GatedStallD),
					.FetchBuffer(FetchBuffer),
					.CacheBusAck(ICacheBusAck),
					.CacheBusAdr(ICacheBusAdr),
					.CacheStall(ICacheStallF),
					.CacheBusRW(CacheBusRW),
					.ReadDataWord(ICacheInstrF),
					.SelHPTW(sv2v_uu_icache_ext_SelHPTW_0),
					.CacheMiss(ICacheMiss),
					.CacheAccess(ICacheAccess),
					.ByteMask(sv2v_uu_icache_ext_ByteMask_0),
					.BeatCount(sv2v_uu_icache_ext_BeatCount_0),
					.SelBusBeat(sv2v_uu_icache_ext_SelBusBeat_0),
					.WriteData(sv2v_uu_icache_ext_WriteData_0),
					.CacheRW(CacheRWF),
					.FlushCache(sv2v_uu_icache_ext_FlushCache_0),
					.NextSet(PCSpillNextF[11:0]),
					.PAdr(PCPF),
					.CacheCommitted(CacheCommittedF),
					.InvalidateCache(InvalidateICacheM),
					.CMOpM(sv2v_uu_icache_ext_CMOpM_0)
				);
				localparam [4216:0] sv2v_uu_ahbcacheinterface_P = P;
				localparam [$signed(sv2v_uu_ahbcacheinterface_P[383-:32]) - 1:0] sv2v_uu_ahbcacheinterface_ext_WriteDataM_0 = 1'sb0;
				localparam [0:0] sv2v_uu_ahbcacheinterface_ext_BusAtomic_0 = 1'sb0;
				localparam [$signed(sv2v_uu_ahbcacheinterface_P[383-:32]) - 1:0] sv2v_uu_ahbcacheinterface_ext_CacheReadDataWordM_0 = 1'sb0;
				ahbcacheinterface #(
					.P(P),
					.BEATSPERLINE(BEATSPERLINE),
					.AHBWLOGBWPL(AHBWLOGBWPL),
					.LINELEN(LINELEN),
					.LLENPOVERAHBW(LLENPOVERAHBW),
					.READ_ONLY_CACHE(1)
				) ahbcacheinterface(
					.HCLK(clk),
					.HRESETn(~reset),
					.HRDATA(HRDATA),
					.Flush(FlushD),
					.CacheBusRW(CacheBusRW),
					.BusCMOZero(1'b0),
					.HSIZE(IFUHSIZE),
					.HBURST(IFUHBURST),
					.HTRANS(IFUHTRANS),
					.HWSTRB(),
					.Funct3(3'b010),
					.HADDR(IFUHADDR),
					.HREADY(IFUHREADY),
					.HWRITE(IFUHWRITE),
					.CacheBusAdr(ICacheBusAdr),
					.BeatCount(),
					.Cacheable(CacheableF),
					.SelBusBeat(),
					.WriteDataM(sv2v_uu_ahbcacheinterface_ext_WriteDataM_0),
					.BusAtomic(sv2v_uu_ahbcacheinterface_ext_BusAtomic_0),
					.CacheBusAck(ICacheBusAck),
					.HWDATA(),
					.CacheableOrFlushCacheM(1'b0),
					.CacheReadDataWordM(sv2v_uu_ahbcacheinterface_ext_CacheReadDataWordM_0),
					.FetchBuffer(FetchBuffer),
					.PAdr(PCPF),
					.BusRW(BusRW),
					.Stall(GatedStallD),
					.BusStall(BusStall),
					.BusCommitted(BusCommittedF)
				);
				mux3 #(.WIDTH(32)) UnCachedDataMux(
					.d0(ICacheInstrF),
					.d1(ShiftUncachedInstr),
					.d2(IROMInstrF),
					.s({SelIROM, ~CacheableF}),
					.y(InstrRawF[31:0])
				);
			end
			else begin : passthrough
				assign IFUHADDR = PCPF;
				wire [1:0] BusRW;
				assign BusRW = (~ITLBMissF & ~SelIROM ? IFURWF : 0);
				assign IFUHSIZE = 3'b010;
				localparam [0:0] sv2v_uu_ahbinterface_ext_BusAtomic_0 = 1'sb0;
				localparam sv2v_uu_ahbinterface_XLEN = $signed(P[4216-:32]);
				localparam [sv2v_uu_ahbinterface_XLEN - 1:0] sv2v_uu_ahbinterface_ext_WriteData_0 = 1'sb0;
				ahbinterface #(
					.XLEN($signed(P[4216-:32])),
					.LSU(1'b0)
				) ahbinterface(
					.HCLK(clk),
					.Flush(FlushD),
					.HRESETn(~reset),
					.HREADY(IFUHREADY),
					.HRDATA(HRDATA),
					.HTRANS(IFUHTRANS),
					.HWRITE(IFUHWRITE),
					.HWDATA(),
					.HWSTRB(),
					.BusRW(BusRW),
					.BusAtomic(sv2v_uu_ahbinterface_ext_BusAtomic_0),
					.ByteMask(),
					.WriteData(sv2v_uu_ahbinterface_ext_WriteData_0),
					.Stall(GatedStallD),
					.BusStall(BusStall),
					.BusCommitted(BusCommittedF),
					.FetchBuffer(FetchBuffer)
				);
				assign CacheCommittedF = 1'sb0;
				if (P[3471]) begin : genblk1
					mux2 #(.WIDTH(32)) UnCachedDataMux2(
						.d0(ShiftUncachedInstr),
						.d1(IROMInstrF),
						.s(SelIROM),
						.y(InstrRawF)
					);
				end
				else begin : genblk1
					assign InstrRawF = ShiftUncachedInstr;
				end
				assign IFUHBURST = 3'b000;
				assign {ICacheMiss, ICacheAccess, ICacheStallF} = 1'sb0;
			end
			if ($signed(P[4216-:32]) == 64) begin : genblk2
				mux4 #(.WIDTH(32)) UncachedShiftInstrMux(
					.d0(FetchBuffer[31:0]),
					.d1(FetchBuffer[47:16]),
					.d2(FetchBuffer[63:32]),
					.d3({16'b0000000000000000, FetchBuffer[63:48]}),
					.s(PCSpillF[2:1]),
					.y(ShiftUncachedInstr)
				);
			end
			else begin : genblk2
				mux2 #(.WIDTH(32)) UncachedShiftInstrMux(
					.d0(FetchBuffer[31:0]),
					.d1({16'b0000000000000000, FetchBuffer[31:16]}),
					.s(PCSpillF[1]),
					.y(ShiftUncachedInstr)
				);
			end
		end
		else begin : nobus
			assign {IFUHADDR, IFUHWRITE, IFUHSIZE, IFUHBURST, IFUHTRANS, BusStall, CacheCommittedF, BusCommittedF, FetchBuffer} = 1'sb0;
			assign {ICacheStallF, ICacheMiss, ICacheAccess} = 1'sb0;
			assign InstrRawF = IROMInstrF;
		end
	endgenerate
	assign IFUCacheBusStallF = ICacheStallF | BusStall;
	assign IFUStallF = IFUCacheBusStallF | SelSpillNextF;
	assign GatedStallD = StallD & ~SelSpillNextF;
	flopenl #(.WIDTH(32)) AlignedInstrRawDFlop(
		.clk(clk),
		.load(reset | FlushD),
		.en(~StallD),
		.d(PostSpillInstrRawF),
		.val(nop),
		.q(InstrRawD)
	);
	generate
		if (P[4086] | P[4085]) begin : genblk5
			mux2 #(.WIDTH($signed(P[4216-:32]))) pcmux2(
				.d0(PC1NextF),
				.d1(NextValidPCE),
				.s(CSRWriteFenceM),
				.y(PC2NextF)
			);
		end
		else begin : genblk5
			assign PC2NextF = PC1NextF;
		end
	endgenerate
	mux3 #(.WIDTH($signed(P[4216-:32]))) pcmux3(
		.d0(PC2NextF),
		.d1(EPCM),
		.d2(TrapVectorM),
		.s({TrapM, RetM}),
		.y(UnalignedPCNextF)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) pcresetmux(
		.d0({UnalignedPCNextF[$signed(P[4216-:32]) - 1:1], 1'b0}),
		.d1(P[$signed(P[4216-:32]) + 3632:3633]),
		.s(reset),
		.y(PCNextF)
	);
	flopen #(.WIDTH($signed(P[4216-:32]))) pcreg(
		.clk(clk),
		.en(~StallF | reset),
		.d(PCNextF),
		.q(PCF)
	);
	assign PCPlus4F = PCF[$signed(P[4216-:32]) - 1:2] + 1;
	generate
		if (P[1754]) begin : pcadd
			always @(*) begin
				if (_sv2v_0)
					;
				if (CompressedF) begin
					if (PCF[1])
						PCPlus2or4F = {PCPlus4F, 2'b00};
					else
						PCPlus2or4F = {PCF[$signed(P[4216-:32]) - 1:2], 2'b10};
				end
				else
					PCPlus2or4F = {PCPlus4F, PCF[1:0]};
			end
		end
		else begin : pcadd
			wire [$signed(P[4216-:32]):1] sv2v_tmp_02717;
			assign sv2v_tmp_02717 = {PCPlus4F, PCF[1:0]};
			always @(*) PCPlus2or4F = sv2v_tmp_02717;
		end
		if (P[1984]) begin : bpred
			bpred #(.P(P)) bpred(
				.clk(clk),
				.reset(reset),
				.StallF(StallF),
				.StallD(StallD),
				.StallE(StallE),
				.StallM(StallM),
				.StallW(StallW),
				.FlushD(FlushD),
				.FlushE(FlushE),
				.FlushM(FlushM),
				.FlushW(FlushW),
				.InstrValidD(InstrValidD),
				.InstrValidE(InstrValidE),
				.BranchD(BranchD),
				.BranchE(BranchE),
				.JumpD(JumpD),
				.JumpE(JumpE),
				.InstrD(InstrD),
				.PCNextF(PCNextF),
				.PCPlus2or4F(PCPlus2or4F),
				.PC1NextF(PC1NextF),
				.PCE(PCE),
				.PCM(PCM),
				.PCSrcE(PCSrcE),
				.IEUAdrE(IEUAdrE),
				.IEUAdrM(IEUAdrM),
				.PCF(PCF),
				.NextValidPCE(NextValidPCE),
				.PCD(PCD),
				.PCLinkE(PCLinkE),
				.IClassM(IClassM),
				.BPWrongE(BPWrongE),
				.PostSpillInstrRawF(PostSpillInstrRawF),
				.BPWrongM(BPWrongM),
				.BPDirWrongM(BPDirWrongM),
				.BTAWrongM(BTAWrongM),
				.RASPredPCWrongM(RASPredPCWrongM),
				.IClassWrongM(IClassWrongM)
			);
		end
		else begin : bpred
			mux2 #(.WIDTH($signed(P[4216-:32]))) pcmux1(
				.d0(PCPlus2or4F),
				.d1(IEUAdrE),
				.s(PCSrcE),
				.y(PC1NextF)
			);
			wire BranchM;
			wire JumpM;
			wire BranchW;
			wire JumpW;
			wire CallD;
			wire CallE;
			wire CallM;
			wire CallW;
			wire ReturnD;
			wire ReturnE;
			wire ReturnM;
			wire ReturnW;
			assign BPWrongE = PCSrcE;
			icpred #(
				.P(P),
				.INSTR_CLASS_PRED(0)
			) icpred(
				.clk(clk),
				.reset(reset),
				.StallD(StallD),
				.StallE(StallE),
				.StallM(StallM),
				.StallW(StallW),
				.FlushD(FlushD),
				.FlushE(FlushE),
				.FlushM(FlushM),
				.PostSpillInstrRawF(PostSpillInstrRawF),
				.InstrD(InstrD),
				.BranchD(BranchD),
				.BranchE(BranchE),
				.JumpD(JumpD),
				.JumpE(JumpE),
				.BranchM(BranchM),
				.BranchW(BranchW),
				.JumpM(JumpM),
				.JumpW(JumpW),
				.CallD(CallD),
				.CallE(CallE),
				.CallM(CallM),
				.CallW(CallW),
				.ReturnD(ReturnD),
				.ReturnE(ReturnE),
				.ReturnM(ReturnM),
				.ReturnW(ReturnW),
				.BTBCallF(1'b0),
				.BTBReturnF(1'b0),
				.BTBJumpF(1'b0),
				.BTBBranchF(1'b0),
				.BPCallF(),
				.BPReturnF(),
				.BPJumpF(),
				.BPBranchF(),
				.IClassWrongM(IClassWrongM),
				.BPReturnWrongD()
			);
			flopenrc #(.WIDTH(1)) PCSrcMReg(
				.clk(clk),
				.reset(reset),
				.clear(FlushM),
				.en(~StallM),
				.d(PCSrcE),
				.q(BPWrongM)
			);
			assign RASPredPCWrongM = 1'b0;
			assign BPDirWrongM = BPWrongM;
			assign BTAWrongM = BPWrongM;
			assign IClassM = {CallM, ReturnM, JumpM, BranchM};
			assign NextValidPCE = PCE;
		end
	endgenerate
	flopenrc #(.WIDTH($signed(P[4216-:32]))) PCDReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallD),
		.d(PCF),
		.q(PCD)
	);
	generate
		if (P[1754]) begin : decomp
			wire IllegalCompInstrD;
			decompress #(.P(P)) decomp(
				.InstrRawD(InstrRawD),
				.InstrD(InstrD),
				.IllegalCompInstrD(IllegalCompInstrD)
			);
			assign IllegalIEUInstrD = IllegalBaseInstrD | IllegalCompInstrD;
		end
		else begin : decomp
			assign InstrD = InstrRawD;
			assign IllegalIEUInstrD = IllegalBaseInstrD;
		end
	endgenerate
	assign IllegalIEUFPUInstrD = IllegalIEUInstrD & (IllegalFPUInstrD | !P[1491]);
	assign BranchMisalignedFaultE = (IEUAdrE[1] & ~P[1754]) & PCSrcE;
	flopenr #(.WIDTH(1)) InstrMisalignedReg(
		.clk(clk),
		.reset(reset),
		.en(~StallM),
		.d(BranchMisalignedFaultE),
		.q(InstrMisalignedFaultM)
	);
	mux2 #(.WIDTH(32)) FlushInstrEMux(
		.d0(InstrD),
		.d1(nop),
		.s(FlushE),
		.y(NextInstrD)
	);
	flopenr #(.WIDTH(32)) InstrEReg(
		.clk(clk),
		.reset(reset),
		.en(~StallE),
		.d(NextInstrD),
		.q(InstrE)
	);
	flopenr #(.WIDTH($signed(P[4216-:32]))) PCEReg(
		.clk(clk),
		.reset(reset),
		.en(~StallE),
		.d(PCD),
		.q(PCE)
	);
	generate
		if ((P[4086] | P[4054]) | P[4053]) begin : genblk9
			mux2 #(.WIDTH(32)) FlushInstrMMux(
				.d0(InstrE),
				.d1(nop),
				.s(FlushM),
				.y(NextInstrE)
			);
			flopenr #(.WIDTH(32)) InstrMReg(
				.clk(clk),
				.reset(reset),
				.en(~StallM),
				.d(NextInstrE),
				.q(InstrM)
			);
		end
		else begin : genblk9
			assign InstrM = 1'sb0;
		end
		if (P[4086] | P[1984]) begin : genblk10
			flopenr #(.WIDTH($signed(P[4216-:32]))) PCMReg(
				.clk(clk),
				.reset(reset),
				.en(~StallM),
				.d(PCE),
				.q(PCM)
			);
		end
		else begin : genblk10
			assign PCM = 1'sb0;
		end
		if (P[1754]) begin : genblk11
			wire CompressedD;
			flopenrc #(.WIDTH(1)) CompressedDReg(
				.clk(clk),
				.reset(reset),
				.clear(FlushD),
				.en(~StallD),
				.d(CompressedF),
				.q(CompressedD)
			);
			flopenrc #(.WIDTH(1)) CompressedEReg(
				.clk(clk),
				.reset(reset),
				.clear(FlushE),
				.en(~StallE),
				.d(CompressedD),
				.q(CompressedE)
			);
			assign PCLinkE = PCE + (CompressedE ? 'd2 : 'd4);
		end
		else begin : genblk11
			assign CompressedE = 1'b0;
			assign PCLinkE = PCE + 'd4;
		end
		if ((P[4086] & P[1754]) | 1) begin : genblk12
			wire CompressedM;
			flopenrc #(.WIDTH(16)) InstrRawEReg(
				.clk(clk),
				.reset(reset),
				.clear(FlushE),
				.en(~StallE),
				.d(InstrRawD[15:0]),
				.q(InstrRawE)
			);
			flopenrc #(.WIDTH(16)) InstrRawMReg(
				.clk(clk),
				.reset(reset),
				.clear(FlushM),
				.en(~StallM),
				.d(InstrRawE),
				.q(InstrRawM)
			);
			flopenrc #(.WIDTH(1)) CompressedMReg(
				.clk(clk),
				.reset(reset),
				.clear(FlushM),
				.en(~StallM),
				.d(CompressedE),
				.q(CompressedM)
			);
			mux2 #(.WIDTH(32)) InstrOrigMux(
				.d0(InstrM),
				.d1({16'b0000000000000000, InstrRawM}),
				.s(CompressedM),
				.y(InstrOrigM)
			);
		end
		else begin : genblk12
			assign InstrOrigM = InstrM;
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module irom (
	clk,
	ce,
	Adr,
	IROMInstrF
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire ce;
	input wire [$signed(P[4216-:32]) - 1:0] Adr;
	output wire [31:0] IROMInstrF;
	localparam XLENBYTES = {{$signed(P[1640-:32]) - 32 {1'b0}}, $signed(P[4216-:32]) / 8};
	localparam ADDR_WDITH = $clog2(P[3342 + $signed(P[1640-:32]):3343] / XLENBYTES);
	localparam OFFSET = $clog2(XLENBYTES);
	wire [$signed(P[4216-:32]) - 1:0] IROMInstrFFull;
	wire [31:0] RawIROMInstrF;
	wire [2:1] AdrD;
	rom1p1r #(
		.ADDR_WIDTH(ADDR_WDITH),
		.DATA_WIDTH($signed(P[4216-:32])),
		.PRELOAD_ENABLED(1)
	) rom(
		.clk(clk),
		.ce(ce),
		.addr(Adr[(ADDR_WDITH + OFFSET) - 1:OFFSET]),
		.dout(IROMInstrFFull)
	);
	generate
		if ($signed(P[4216-:32]) == 32) begin : genblk1
			assign RawIROMInstrF = IROMInstrFFull;
		end
		else begin : genblk1
			flopen #(.WIDTH(1)) AdrReg2(
				.clk(clk),
				.en(ce),
				.d(Adr[2]),
				.q(AdrD[2])
			);
			assign RawIROMInstrF = (AdrD[2] ? IROMInstrFFull[63:32] : IROMInstrFFull[31:0]);
		end
		if (P[1754]) begin : genblk2
			flopen #(.WIDTH(1)) AdrReg1(
				.clk(clk),
				.en(ce),
				.d(Adr[1]),
				.q(AdrD[1])
			);
			assign IROMInstrF = (AdrD[1] ? {16'b0000000000000000, RawIROMInstrF[31:16]} : RawIROMInstrF);
		end
		else begin : genblk2
			assign IROMInstrF = RawIROMInstrF;
		end
	endgenerate
endmodule
module spill (
	clk,
	reset,
	StallF,
	FlushD,
	PCF,
	PCPlus4F,
	PCNextF,
	InstrRawF,
	IFUCacheBusStallF,
	ITLBMissOrUpdateAF,
	CacheableF,
	PCSpillNextF,
	PCSpillF,
	SelSpillNextF,
	PostSpillInstrRawF,
	CompressedF
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallF;
	input wire FlushD;
	input wire [$signed(P[4216-:32]) - 1:0] PCF;
	input wire [$signed(P[4216-:32]) - 1:2] PCPlus4F;
	input wire [$signed(P[4216-:32]) - 1:0] PCNextF;
	input wire [31:0] InstrRawF;
	input wire IFUCacheBusStallF;
	input wire ITLBMissOrUpdateAF;
	input wire CacheableF;
	output wire [$signed(P[4216-:32]) - 1:0] PCSpillNextF;
	output wire [$signed(P[4216-:32]) - 1:0] PCSpillF;
	output wire SelSpillNextF;
	output wire [31:0] PostSpillInstrRawF;
	output reg CompressedF;
	reg [1:0] CurrState;
	reg [1:0] NextState;
	wire [$signed(P[4216-:32]) - 1:0] PCPlus2NextF;
	wire [$signed(P[4216-:32]) - 1:0] PCPlus2F;
	wire TakeSpillF;
	wire SpillF;
	wire SelSpillF;
	wire SpillSaveF;
	wire [15:0] InstrFirstHalfF;
	wire EarlyCompressedF;
	mux2 #(.WIDTH($signed(P[4216-:32]))) pcplus2mux(
		.d0({PCF[$signed(P[4216-:32]) - 1:2], 2'b10}),
		.d1({PCPlus4F, 2'b00}),
		.s(PCF[1]),
		.y(PCPlus2NextF)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) pcnextspillmux(
		.d0(PCNextF),
		.d1(PCPlus2NextF),
		.s(SelSpillNextF & ~FlushD),
		.y(PCSpillNextF)
	);
	flopr #(.WIDTH($signed(P[4216-:32]))) pcplus2reg(
		.clk(clk),
		.reset(reset),
		.d(PCPlus2NextF),
		.q(PCPlus2F)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) pcspillmux(
		.d0(PCF),
		.d1(PCPlus2F),
		.s(SelSpillF),
		.y(PCSpillF)
	);
	generate
		if (P[4050]) begin : genblk1
			wire SpillCachedF;
			wire SpillUncachedF;
			assign SpillCachedF = &PCF[$clog2($signed(P[3825-:32]) / 32) + 1:1];
			assign SpillUncachedF = PCF[1];
			assign SpillF = (CacheableF ? SpillCachedF : SpillUncachedF);
		end
		else begin : genblk1
			assign SpillF = PCF[1];
		end
	endgenerate
	assign TakeSpillF = ((SpillF & ~EarlyCompressedF) & ~IFUCacheBusStallF) & ~ITLBMissOrUpdateAF;
	always @(posedge clk)
		if (reset | FlushD)
			CurrState <= 2'd0;
		else
			CurrState <= NextState;
	always @(*) begin
		if (_sv2v_0)
			;
		case (CurrState)
			2'd0:
				if (TakeSpillF)
					NextState = 2'd1;
				else
					NextState = 2'd0;
			2'd1:
				if (StallF)
					NextState = 2'd1;
				else
					NextState = 2'd0;
			default: NextState = 2'd0;
		endcase
	end
	assign SelSpillF = CurrState == 2'd1;
	assign SelSpillNextF = ((CurrState == 2'd0) & TakeSpillF) | ((CurrState == 2'd1) & IFUCacheBusStallF);
	assign SpillSaveF = ((CurrState == 2'd0) & TakeSpillF) & ~FlushD;
	flopenr #(.WIDTH(16)) SpillInstrReg(
		.clk(clk),
		.reset(reset),
		.en(SpillSaveF),
		.d(InstrRawF[15:0]),
		.q(InstrFirstHalfF)
	);
	mux2 #(.WIDTH(32)) postspillmux(
		.d0(InstrRawF),
		.d1({InstrRawF[15:0], InstrFirstHalfF}),
		.s(SelSpillF),
		.y(PostSpillInstrRawF)
	);
	always @(*) begin
		if (_sv2v_0)
			;
		if (PostSpillInstrRawF[1:0] != 2'b11)
			CompressedF = 1'b1;
		else
			CompressedF = 1'b0;
	end
	assign EarlyCompressedF = ~(&InstrRawF[1:0]);
	initial _sv2v_0 = 0;
endmodule
module align (
	clk,
	reset,
	StallM,
	FlushM,
	IEUAdrM,
	IEUAdrE,
	Funct3M,
	FpLoadStoreM,
	MemRWM,
	DCacheReadDataWordM,
	CacheBusHPWTStall,
	SelHPTW,
	ByteMaskM,
	ByteMaskExtendedM,
	LSUWriteDataM,
	ByteMaskSpillM,
	LSUWriteDataSpillM,
	IEUAdrSpillE,
	IEUAdrSpillM,
	IEUAdrxTvalM,
	SelSpillE,
	DCacheReadDataWordSpillM,
	SpillStallM
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallM;
	input wire FlushM;
	input wire [$signed(P[4216-:32]) - 1:0] IEUAdrM;
	input wire [$signed(P[4216-:32]) - 1:0] IEUAdrE;
	input wire [2:0] Funct3M;
	input wire FpLoadStoreM;
	input wire [1:0] MemRWM;
	input wire [($signed(P[383-:32]) * 2) - 1:0] DCacheReadDataWordM;
	input wire CacheBusHPWTStall;
	input wire SelHPTW;
	input wire [($signed(P[383-:32]) - 1) / 8:0] ByteMaskM;
	input wire [($signed(P[383-:32]) - 1) / 8:0] ByteMaskExtendedM;
	input wire [$signed(P[383-:32]) - 1:0] LSUWriteDataM;
	output wire [(($signed(P[383-:32]) * 2) - 1) / 8:0] ByteMaskSpillM;
	output wire [($signed(P[383-:32]) * 2) - 1:0] LSUWriteDataSpillM;
	output wire [$signed(P[4216-:32]) - 1:0] IEUAdrSpillE;
	output wire [$signed(P[4216-:32]) - 1:0] IEUAdrSpillM;
	output wire [$signed(P[4216-:32]) - 1:0] IEUAdrxTvalM;
	output wire SelSpillE;
	output wire [$signed(P[383-:32]) - 1:0] DCacheReadDataWordSpillM;
	output wire SpillStallM;
	localparam LLENINBYTES = $signed(P[383-:32]) / 8;
	localparam OFFSET_BIT_POS = $clog2($signed(P[3921-:32]) / 8);
	reg [1:0] CurrState;
	reg [1:0] NextState;
	wire ValidSpillM;
	wire SelSpillM;
	wire SpillSaveM;
	wire [$signed(P[383-:32]) - 1:0] ReadDataWordFirstHalfM;
	wire MisalignedM;
	wire [($signed(P[383-:32]) * 2) - 1:0] ReadDataWordSpillAllM;
	wire [($signed(P[383-:32]) * 2) - 1:0] ReadDataWordSpillShiftedM;
	wire [$signed(P[4216-:32]) - 1:0] IEUAdrIncrementM;
	localparam OFFSET_LEN = $clog2(LLENINBYTES);
	reg [$clog2(LLENINBYTES) - 1:0] AccessByteOffsetM;
	wire [$clog2(LLENINBYTES) + 2:0] ShiftAmount;
	reg PotentialSpillM;
	wire [($signed(P[383-:32]) * 3) - 1:0] LSUWriteDataShiftedExtM;
	assign IEUAdrIncrementM = IEUAdrM + LLENINBYTES;
	mux2 #(.WIDTH($signed(P[4216-:32]))) ieuadrspillemux(
		.d0(IEUAdrE),
		.d1(IEUAdrIncrementM),
		.s(SelSpillE),
		.y(IEUAdrSpillE)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) ieuadrspillmmux(
		.d0(IEUAdrM),
		.d1(IEUAdrIncrementM),
		.s(SelSpillM),
		.y(IEUAdrSpillM)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) ieuadrxtvalmmux(
		.d0(IEUAdrM),
		.d1({IEUAdrIncrementM[$signed(P[4216-:32]) - 1:OFFSET_LEN], {{OFFSET_LEN} {1'b0}}}),
		.s(SelSpillM),
		.y(IEUAdrxTvalM)
	);
	always @(*) begin
		if (_sv2v_0)
			;
		case (Funct3M & {FpLoadStoreM, 2'b11})
			3'b000: AccessByteOffsetM = 1'sb0;
			3'b001: AccessByteOffsetM = {{OFFSET_LEN - 1 {1'b0}}, IEUAdrM[0]};
			3'b010: AccessByteOffsetM = {{OFFSET_LEN - 2 {1'b0}}, IEUAdrM[1:0]};
			3'b011:
				if ($signed(P[383-:32]) >= 64)
					AccessByteOffsetM = {{OFFSET_LEN - 3 {1'b0}}, IEUAdrM[2:0]};
				else
					AccessByteOffsetM = 1'sb0;
			3'b100:
				if ($signed(P[383-:32]) == 128)
					AccessByteOffsetM = IEUAdrM[OFFSET_LEN - 1:0];
				else
					AccessByteOffsetM = IEUAdrM[OFFSET_LEN - 1:0];
			default: AccessByteOffsetM = 1'sb0;
		endcase
		case (Funct3M[1:0])
			2'b00: PotentialSpillM = 1'b0;
			2'b01: PotentialSpillM = IEUAdrM[OFFSET_BIT_POS - 1:1] == {((OFFSET_BIT_POS - 1) >= 1 ? OFFSET_BIT_POS - 1 : 3 - OFFSET_BIT_POS) * 1 {1'sb1}};
			2'b10: PotentialSpillM = IEUAdrM[OFFSET_BIT_POS - 1:2] == {((OFFSET_BIT_POS - 1) >= 2 ? OFFSET_BIT_POS - 2 : 4 - OFFSET_BIT_POS) * 1 {1'sb1}};
			2'b11: PotentialSpillM = IEUAdrM[OFFSET_BIT_POS - 1:3] == {((OFFSET_BIT_POS - 1) >= 3 ? OFFSET_BIT_POS - 3 : 5 - OFFSET_BIT_POS) * 1 {1'sb1}};
			default: PotentialSpillM = 1'b0;
		endcase
	end
	assign MisalignedM = |MemRWM & (AccessByteOffsetM != 0);
	assign ValidSpillM = (MisalignedM & PotentialSpillM) & ~CacheBusHPWTStall;
	always @(posedge clk)
		if (reset | FlushM)
			CurrState <= 2'd0;
		else
			CurrState <= NextState;
	always @(*) begin
		if (_sv2v_0)
			;
		case (CurrState)
			2'd0:
				if (ValidSpillM)
					NextState = 2'd1;
				else
					NextState = 2'd0;
			2'd1:
				if (StallM)
					NextState = 2'd1;
				else
					NextState = 2'd0;
			default: NextState = 2'd0;
		endcase
	end
	assign SelSpillM = CurrState == 2'd1;
	assign SelSpillE = ((CurrState == 2'd0) & ValidSpillM) | ((CurrState == 2'd1) & CacheBusHPWTStall);
	assign SpillSaveM = ((CurrState == 2'd0) & ValidSpillM) & ~FlushM;
	assign SpillStallM = SelSpillE;
	flopenr #(.WIDTH($signed(P[383-:32]))) SpillDataReg(
		.clk(clk),
		.reset(reset),
		.en(SpillSaveM),
		.d(DCacheReadDataWordM[$signed(P[383-:32]) - 1:0]),
		.q(ReadDataWordFirstHalfM)
	);
	mux2 #(.WIDTH(2 * $signed(P[383-:32]))) postspillmux(
		.d0(DCacheReadDataWordM),
		.d1({DCacheReadDataWordM[$signed(P[383-:32]) - 1:0], ReadDataWordFirstHalfM}),
		.s(SelSpillM & ~SelHPTW),
		.y(ReadDataWordSpillAllM)
	);
	assign ShiftAmount = (SelHPTW ? {(($clog2(LLENINBYTES) + 2) >= 0 ? $clog2(LLENINBYTES) + 3 : 1 - ($clog2(LLENINBYTES) + 2)) {1'sb0}} : {AccessByteOffsetM, 3'b000});
	assign ReadDataWordSpillShiftedM = ReadDataWordSpillAllM >> ShiftAmount;
	assign DCacheReadDataWordSpillM = ReadDataWordSpillShiftedM[$signed(P[383-:32]) - 1:0];
	assign LSUWriteDataShiftedExtM = {LSUWriteDataM, LSUWriteDataM, LSUWriteDataM} << ShiftAmount;
	assign LSUWriteDataSpillM = LSUWriteDataShiftedExtM[($signed(P[383-:32]) * 3) - 1:$signed(P[383-:32])];
	mux3 #(.WIDTH((2 * $signed(P[383-:32])) / 8)) bytemaskspillmux(
		.d0({ByteMaskExtendedM, ByteMaskM}),
		.d1({{{$signed(P[383-:32]) / 8} {1'b0}}, ByteMaskM}),
		.d2({{{$signed(P[383-:32]) / 8} {1'b0}}, ByteMaskExtendedM}),
		.s({SelSpillM, SelSpillE}),
		.y(ByteMaskSpillM)
	);
	initial _sv2v_0 = 0;
endmodule
module amoalu (
	ReadDataM,
	IHWriteDataM,
	LSUFunct7M,
	LSUFunct3M,
	AMOResultM
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[4216-:32]) - 1:0] ReadDataM;
	input wire [$signed(P[4216-:32]) - 1:0] IHWriteDataM;
	input wire [6:0] LSUFunct7M;
	input wire [2:0] LSUFunct3M;
	output reg [$signed(P[4216-:32]) - 1:0] AMOResultM;
	wire [$signed(P[4216-:32]) - 1:0] a;
	wire [$signed(P[4216-:32]) - 1:0] b;
	reg [$signed(P[4216-:32]) - 1:0] y;
	wire lt;
	wire cmp;
	wire sngd;
	wire sngd32;
	wire eq32;
	wire lt32;
	wire w64;
	assign a = ReadDataM;
	assign b = IHWriteDataM;
	assign sngd = ~LSUFunct7M[5];
	assign w64 = LSUFunct3M[1:0] == 2'b10;
	assign sngd32 = sngd & (($signed(P[4216-:32]) == 32) | w64);
	comparator #(.WIDTH(32)) cmp32(
		.a(a[31:0]),
		.b(b[31:0]),
		.sgnd(sngd32),
		.flags({eq32, lt32})
	);
	generate
		if ($signed(P[4216-:32]) == 32) begin : genblk1
			assign lt = lt32;
		end
		else begin : genblk1
			wire equpper;
			wire ltupper;
			wire lt64;
			comparator #(.WIDTH(32)) cmpupper(
				.a(a[63:32]),
				.b(b[63:32]),
				.sgnd(sngd),
				.flags({equpper, ltupper})
			);
			assign lt64 = ltupper | (equpper & lt32);
			assign lt = (w64 ? lt32 : lt64);
		end
	endgenerate
	assign cmp = lt ^ LSUFunct7M[4];
	always @(*) begin
		if (_sv2v_0)
			;
		case (LSUFunct7M[6:2])
			5'b00001: y = b;
			5'b00000: y = a + b;
			5'b00100: y = a ^ b;
			5'b01100: y = a & b;
			5'b01000: y = a | b;
			5'b10000: y = (cmp ? a : b);
			5'b10100: y = (cmp ? a : b);
			5'b11000: y = (cmp ? a : b);
			5'b11100: y = (cmp ? a : b);
			default: y = 1'sbx;
		endcase
	end
	generate
		if ($signed(P[4216-:32]) == 32) begin : sext
			wire [$signed(P[4216-:32]):1] sv2v_tmp_250F8;
			assign sv2v_tmp_250F8 = y;
			always @(*) AMOResultM = sv2v_tmp_250F8;
		end
		else begin : sext
			always @(*) begin
				if (_sv2v_0)
					;
				if (w64)
					AMOResultM = {{32 {y[31]}}, y[31:0]};
				else
					AMOResultM = y;
			end
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module atomic (
	clk,
	reset,
	StallW,
	ReadDataM,
	IHWriteDataM,
	PAdrM,
	LSUFunct7M,
	LSUFunct3M,
	LSUAtomicM,
	PreLSURWM,
	LSUFlushW,
	IMAWriteDataM,
	SquashSCW,
	LSURWM
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallW;
	input wire [$signed(P[4216-:32]) - 1:0] ReadDataM;
	input wire [$signed(P[4216-:32]) - 1:0] IHWriteDataM;
	input wire [$signed(P[1640-:32]) - 1:0] PAdrM;
	input wire [6:0] LSUFunct7M;
	input wire [2:0] LSUFunct3M;
	input wire [1:0] LSUAtomicM;
	input wire [1:0] PreLSURWM;
	input wire LSUFlushW;
	output wire [$signed(P[4216-:32]) - 1:0] IMAWriteDataM;
	output wire SquashSCW;
	output wire [1:0] LSURWM;
	wire [$signed(P[4216-:32]) - 1:0] AMOResultM;
	wire MemReadM;
	generate
		if (P[4054]) begin : genblk1
			amoalu #(.P(P)) amoalu(
				.ReadDataM(ReadDataM),
				.IHWriteDataM(IHWriteDataM),
				.LSUFunct7M(LSUFunct7M),
				.LSUFunct3M(LSUFunct3M),
				.AMOResultM(AMOResultM)
			);
			mux2 #(.WIDTH($signed(P[4216-:32]))) wdmux(
				.d0(IHWriteDataM),
				.d1(AMOResultM),
				.s(LSUAtomicM[1]),
				.y(IMAWriteDataM)
			);
		end
		else begin : genblk1
			assign IMAWriteDataM = IHWriteDataM;
		end
		if (P[4053]) begin : genblk2
			assign MemReadM = PreLSURWM[1] & ~LSUFlushW;
			lrsc #(.P(P)) lrsc(
				.clk(clk),
				.reset(reset),
				.StallW(StallW),
				.MemReadM(MemReadM),
				.PreLSURWM(PreLSURWM),
				.LSUAtomicM(LSUAtomicM),
				.PAdrM(PAdrM),
				.SquashSCW(SquashSCW),
				.LSURWM(LSURWM)
			);
		end
		else begin : genblk2
			assign SquashSCW = 0;
			assign LSURWM = PreLSURWM;
		end
	endgenerate
endmodule
module dtim (
	clk,
	reset,
	FlushW,
	ce,
	MemRWM,
	DTIMAdr,
	WriteDataM,
	ByteMaskM,
	ReadDataWordM
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire FlushW;
	input wire ce;
	input wire [1:0] MemRWM;
	input wire [$signed(P[1640-:32]) - 1:0] DTIMAdr;
	input wire [$signed(P[383-:32]) - 1:0] WriteDataM;
	input wire [($signed(P[383-:32]) / 8) - 1:0] ByteMaskM;
	output wire [$signed(P[383-:32]) - 1:0] ReadDataWordM;
	wire we;
	localparam LLENBYTES = $signed(P[383-:32]) / 8;
	localparam DEPTH = P[3535-:64] / LLENBYTES;
	localparam ADDR_WDITH = $clog2(DEPTH);
	localparam OFFSET = $clog2(LLENBYTES);
	assign we = MemRWM[0] & ~FlushW;
	ram1p1rwbe #(
		.USE_SRAM(P[1743]),
		.DEPTH(DEPTH),
		.WIDTH($signed(P[383-:32]))
	) ram(
		.clk(clk),
		.ce(ce),
		.we(we),
		.bwe(ByteMaskM),
		.addr(DTIMAdr[(ADDR_WDITH + OFFSET) - 1:OFFSET]),
		.dout(ReadDataWordM),
		.din(WriteDataM)
	);
endmodule
module endianswap (
	BigEndianM,
	a,
	y
);
	reg _sv2v_0;
	parameter LEN = 0;
	input wire BigEndianM;
	input wire [LEN - 1:0] a;
	output reg [LEN - 1:0] y;
	generate
		if (LEN == 128) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				if (BigEndianM) begin
					y[127:120] = a[7:0];
					y[119:112] = a[15:8];
					y[111:104] = a[23:16];
					y[103:96] = a[31:24];
					y[95:88] = a[39:32];
					y[87:80] = a[47:40];
					y[79:72] = a[55:48];
					y[71:64] = a[63:56];
					y[63:56] = a[71:64];
					y[55:48] = a[79:72];
					y[47:40] = a[87:80];
					y[39:32] = a[95:88];
					y[31:24] = a[103:96];
					y[23:16] = a[111:104];
					y[15:8] = a[119:112];
					y[7:0] = a[127:120];
				end
				else
					y = a;
			end
		end
		else if (LEN == 64) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				if (BigEndianM) begin
					y[63:56] = a[7:0];
					y[55:48] = a[15:8];
					y[47:40] = a[23:16];
					y[39:32] = a[31:24];
					y[31:24] = a[39:32];
					y[23:16] = a[47:40];
					y[15:8] = a[55:48];
					y[7:0] = a[63:56];
				end
				else
					y = a;
			end
		end
		else begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				if (BigEndianM) begin
					y[31:24] = a[7:0];
					y[23:16] = a[15:8];
					y[15:8] = a[23:16];
					y[7:0] = a[31:24];
				end
				else
					y = a;
			end
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module lrsc (
	clk,
	reset,
	StallW,
	MemReadM,
	PreLSURWM,
	LSURWM,
	LSUAtomicM,
	PAdrM,
	SquashSCW
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallW;
	input wire MemReadM;
	input wire [1:0] PreLSURWM;
	output wire [1:0] LSURWM;
	input wire [1:0] LSUAtomicM;
	input wire [$signed(P[1640-:32]) - 1:0] PAdrM;
	output wire SquashSCW;
	localparam RESERVATION_SET_SIZE_IN_BYTES = $signed(P[4216-:32]) / 8;
	localparam RESERVATION_SET_ADDRESS_BITS = $clog2(RESERVATION_SET_SIZE_IN_BYTES);
	wire [$signed(P[1640-:32]) - 1:RESERVATION_SET_ADDRESS_BITS] ReservationPAdrW;
	reg ReservationValidM;
	wire ReservationValidW;
	wire lrM;
	wire scM;
	wire WriteAdrMatchM;
	wire SquashSCM;
	assign lrM = MemReadM & LSUAtomicM[0];
	assign scM = PreLSURWM[0] & LSUAtomicM[0];
	assign WriteAdrMatchM = (PreLSURWM[0] & (PAdrM[$signed(P[1640-:32]) - 1:RESERVATION_SET_ADDRESS_BITS] == ReservationPAdrW)) & ReservationValidW;
	assign SquashSCM = scM & ~WriteAdrMatchM;
	assign LSURWM = (SquashSCM ? 2'b00 : PreLSURWM);
	always @(*) begin
		if (_sv2v_0)
			;
		if (lrM)
			ReservationValidM = 1'b1;
		else if (scM)
			ReservationValidM = 1'b0;
		else
			ReservationValidM = ReservationValidW;
	end
	flopenr #(.WIDTH($signed(P[1640-:32]) - RESERVATION_SET_ADDRESS_BITS)) resadrreg(
		.clk(clk),
		.reset(reset),
		.en(lrM & ~StallW),
		.d(PAdrM[$signed(P[1640-:32]) - 1:RESERVATION_SET_ADDRESS_BITS]),
		.q(ReservationPAdrW)
	);
	flopenr #(.WIDTH(1)) resvldreg(
		.clk(clk),
		.reset(reset),
		.en(~StallW),
		.d(ReservationValidM),
		.q(ReservationValidW)
	);
	flopenr #(.WIDTH(1)) squashreg(
		.clk(clk),
		.reset(reset),
		.en(~StallW),
		.d(SquashSCM),
		.q(SquashSCW)
	);
	initial _sv2v_0 = 0;
endmodule
module lsu (
	clk,
	reset,
	StallM,
	FlushM,
	StallW,
	FlushW,
	LSUStallM,
	MemRWE,
	MemRWM,
	Funct3M,
	Funct7M,
	AtomicM,
	FlushDCacheM,
	CMOpM,
	LSUPrefetchM,
	CommittedM,
	SquashSCW,
	DCacheMiss,
	DCacheAccess,
	IEUAdrE,
	IEUAdrM,
	WriteDataM,
	ReadDataW,
	PrivilegeModeW,
	BigEndianM,
	sfencevmaM,
	DCacheStallM,
	IEUAdrxTvalM,
	FWriteDataM,
	FpLoadStoreM,
	LoadPageFaultM,
	StoreAmoPageFaultM,
	LoadMisalignedFaultM,
	LoadAccessFaultM,
	HPTWInstrAccessFaultF,
	HPTWInstrPageFaultF,
	StoreAmoMisalignedFaultM,
	StoreAmoAccessFaultM,
	LSUHADDR,
	HRDATA,
	LSUHWDATA,
	LSUHREADY,
	LSUHWRITE,
	LSUHSIZE,
	LSUHBURST,
	LSUHTRANS,
	LSUHWSTRB,
	SATP_REGW,
	STATUS_MXR,
	STATUS_SUM,
	STATUS_MPRV,
	STATUS_MPP,
	ENVCFG_PBMTE,
	ENVCFG_ADUE,
	PCSpillF,
	ITLBMissOrUpdateAF,
	PTE,
	PageType,
	ITLBWriteF,
	SelHPTW,
	PMPCFG_ARRAY_REGW,
	PMPADDR_ARRAY_REGW
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallM;
	input wire FlushM;
	input wire StallW;
	input wire FlushW;
	output wire LSUStallM;
	input wire [1:0] MemRWE;
	input wire [1:0] MemRWM;
	input wire [2:0] Funct3M;
	input wire [6:0] Funct7M;
	input wire [1:0] AtomicM;
	input wire FlushDCacheM;
	input wire [3:0] CMOpM;
	input wire LSUPrefetchM;
	output wire CommittedM;
	output wire SquashSCW;
	output wire DCacheMiss;
	output wire DCacheAccess;
	input wire [$signed(P[4216-:32]) - 1:0] IEUAdrE;
	output wire [$signed(P[4216-:32]) - 1:0] IEUAdrM;
	input wire [$signed(P[4216-:32]) - 1:0] WriteDataM;
	output wire [$signed(P[383-:32]) - 1:0] ReadDataW;
	input wire [1:0] PrivilegeModeW;
	input wire BigEndianM;
	input wire sfencevmaM;
	output wire DCacheStallM;
	output wire [$signed(P[4216-:32]) - 1:0] IEUAdrxTvalM;
	input wire [$signed(P[901-:32]) - 1:0] FWriteDataM;
	input wire FpLoadStoreM;
	output wire LoadPageFaultM;
	output wire StoreAmoPageFaultM;
	output wire LoadMisalignedFaultM;
	output wire LoadAccessFaultM;
	output wire HPTWInstrAccessFaultF;
	output wire HPTWInstrPageFaultF;
	output wire StoreAmoMisalignedFaultM;
	output wire StoreAmoAccessFaultM;
	output wire [$signed(P[1640-:32]) - 1:0] LSUHADDR;
	input wire [$signed(P[4216-:32]) - 1:0] HRDATA;
	output wire [$signed(P[4216-:32]) - 1:0] LSUHWDATA;
	input wire LSUHREADY;
	output wire LSUHWRITE;
	output wire [2:0] LSUHSIZE;
	output wire [2:0] LSUHBURST;
	output wire [1:0] LSUHTRANS;
	output wire [($signed(P[4216-:32]) / 8) - 1:0] LSUHWSTRB;
	input wire [$signed(P[4216-:32]) - 1:0] SATP_REGW;
	input wire STATUS_MXR;
	input wire STATUS_SUM;
	input wire STATUS_MPRV;
	input wire [1:0] STATUS_MPP;
	input wire ENVCFG_PBMTE;
	input wire ENVCFG_ADUE;
	input wire [$signed(P[4216-:32]) - 1:0] PCSpillF;
	input wire ITLBMissOrUpdateAF;
	output wire [$signed(P[4216-:32]) - 1:0] PTE;
	output wire [1:0] PageType;
	output wire ITLBWriteF;
	output wire SelHPTW;
	input wire [($signed(P[3728-:32]) * 8) - 1:0] PMPCFG_ARRAY_REGW;
	input wire [(($signed(P[1640-:32]) - 3) >= 0 ? ($signed(P[3728-:32]) * ($signed(P[1640-:32]) - 2)) - 1 : ($signed(P[3728-:32]) * (4 - $signed(P[1640-:32]))) + ($signed(P[1640-:32]) - 4)):(($signed(P[1640-:32]) - 3) >= 0 ? 0 : $signed(P[1640-:32]) - 3)] PMPADDR_ARRAY_REGW;
	localparam [0:0] MISALIGN_SUPPORT = P[4059] & P[4051];
	localparam MLEN = (MISALIGN_SUPPORT ? 2 * $signed(P[383-:32]) : $signed(P[383-:32]));
	wire [$signed(P[4216-:32]) + 1:0] IEUAdrExtM;
	wire [$signed(P[4216-:32]) + 1:0] IEUAdrExtE;
	wire [$signed(P[1640-:32]) - 1:0] PAdrM;
	wire [$signed(P[4216-:32]) + 1:0] IHAdrM;
	wire [1:0] PreLSURWM;
	wire [1:0] LSURWM;
	wire [2:0] LSUFunct3M;
	wire [6:0] LSUFunct7M;
	wire [1:0] LSUAtomicM;
	wire GatedStallW;
	wire LSUBusStallM;
	wire HPTWStall;
	wire DCacheBusStallM;
	wire CacheBusHPWTStall;
	wire SelSpillE;
	wire CacheableM;
	wire BusCommittedM;
	wire DCacheCommittedM;
	wire [$signed(P[383-:32]) - 1:0] DTIMReadDataWordM;
	wire [MLEN - 1:0] DCacheReadDataWordM;
	wire [MLEN - 1:0] LSUWriteDataSpillM;
	wire [(MLEN / 8) - 1:0] ByteMaskSpillM;
	wire [$signed(P[383-:32]) - 1:0] DCacheReadDataWordSpillM;
	wire [$signed(P[383-:32]) - 1:0] ReadDataWordMuxM;
	wire [$signed(P[383-:32]) - 1:0] LittleEndianReadDataWordM;
	wire [$signed(P[383-:32]) - 1:0] ReadDataM;
	wire [$signed(P[4216-:32]) - 1:0] IHWriteDataM;
	wire [$signed(P[4216-:32]) - 1:0] IMAWriteDataM;
	wire [$signed(P[383-:32]) - 1:0] IMAFWriteDataM;
	wire [$signed(P[383-:32]) - 1:0] LittleEndianWriteDataM;
	wire [$signed(P[383-:32]) - 1:0] LSUWriteDataM;
	wire [($signed(P[383-:32]) - 1) / 8:0] ByteMaskM;
	wire [($signed(P[383-:32]) - 1) / 8:0] ByteMaskExtendedM;
	wire [1:0] MemRWSpillM;
	wire SpillStallM;
	wire DTLBMissM;
	wire DTLBWriteM;
	wire LSULoadAccessFaultM;
	wire LSUStoreAmoAccessFaultM;
	wire HPTWFlushW;
	wire LSUFlushW;
	wire SelDTIM;
	wire [$signed(P[4216-:32]) - 1:0] WriteDataZM;
	wire LSULoadPageFaultM;
	wire LSUStoreAmoPageFaultM;
	wire DTLBMissOrUpdateDAM;
	flopenrc #(.WIDTH($signed(P[4216-:32]))) AddressMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(IEUAdrE),
		.q(IEUAdrM)
	);
	generate
		if (MISALIGN_SUPPORT) begin : ziccslm_align
			wire [$signed(P[4216-:32]) - 1:0] IEUAdrSpillE;
			wire [$signed(P[4216-:32]) - 1:0] IEUAdrSpillM;
			align #(.P(P)) align(
				.clk(clk),
				.reset(reset),
				.StallM(StallM),
				.FlushM(FlushM),
				.IEUAdrE(IEUAdrE),
				.IEUAdrM(IEUAdrM),
				.Funct3M(Funct3M),
				.FpLoadStoreM(FpLoadStoreM),
				.MemRWM(MemRWM),
				.DCacheReadDataWordM(DCacheReadDataWordM),
				.CacheBusHPWTStall(CacheBusHPWTStall),
				.SelHPTW(SelHPTW),
				.ByteMaskM(ByteMaskM),
				.ByteMaskExtendedM(ByteMaskExtendedM),
				.LSUWriteDataM(LSUWriteDataM),
				.ByteMaskSpillM(ByteMaskSpillM),
				.LSUWriteDataSpillM(LSUWriteDataSpillM),
				.IEUAdrSpillE(IEUAdrSpillE),
				.IEUAdrSpillM(IEUAdrSpillM),
				.IEUAdrxTvalM(IEUAdrxTvalM),
				.SelSpillE(SelSpillE),
				.DCacheReadDataWordSpillM(DCacheReadDataWordSpillM),
				.SpillStallM(SpillStallM)
			);
			assign IEUAdrExtM = {2'b00, IEUAdrSpillM};
			assign IEUAdrExtE = {2'b00, IEUAdrSpillE};
		end
		else begin : no_ziccslm_align
			assign IEUAdrExtM = {2'b00, IEUAdrM};
			assign IEUAdrExtE = {2'b00, IEUAdrE};
			assign SelSpillE = 1'b0;
			assign DCacheReadDataWordSpillM = DCacheReadDataWordM;
			assign ByteMaskSpillM = ByteMaskM;
			assign LSUWriteDataSpillM = LSUWriteDataM;
			assign MemRWSpillM = MemRWM;
			assign {SpillStallM} = 1'b0;
			assign IEUAdrxTvalM = IEUAdrM;
		end
		if (P[4061]) begin : cboz
			assign WriteDataZM = (CMOpM[3] ? 0 : WriteDataM);
		end
		else begin : cboz
			assign WriteDataZM = WriteDataM;
		end
		if (P[4067]) begin : hptw
			hptw #(.P(P)) hptw(
				.clk(clk),
				.reset(reset),
				.MemRWM(MemRWM),
				.AtomicM(AtomicM),
				.ITLBMissOrUpdateAF(ITLBMissOrUpdateAF),
				.ITLBWriteF(ITLBWriteF),
				.DTLBMissOrUpdateDAM(DTLBMissOrUpdateDAM),
				.DTLBWriteM(DTLBWriteM),
				.FlushW(FlushW),
				.DCacheBusStallM(DCacheBusStallM),
				.SATP_REGW(SATP_REGW),
				.PCSpillF(PCSpillF),
				.STATUS_MXR(STATUS_MXR),
				.STATUS_SUM(STATUS_SUM),
				.STATUS_MPRV(STATUS_MPRV),
				.STATUS_MPP(STATUS_MPP),
				.ENVCFG_ADUE(ENVCFG_ADUE),
				.PrivilegeModeW(PrivilegeModeW),
				.ReadDataM(ReadDataM[$signed(P[4216-:32]) - 1:0]),
				.WriteDataM(WriteDataZM),
				.Funct3M(Funct3M),
				.LSUFunct3M(LSUFunct3M),
				.Funct7M(Funct7M),
				.LSUFunct7M(LSUFunct7M),
				.IEUAdrExtM(IEUAdrExtM),
				.PTE(PTE),
				.IHWriteDataM(IHWriteDataM),
				.PageType(PageType),
				.PreLSURWM(PreLSURWM),
				.LSUAtomicM(LSUAtomicM),
				.IHAdrM(IHAdrM),
				.HPTWStall(HPTWStall),
				.SelHPTW(SelHPTW),
				.HPTWFlushW(HPTWFlushW),
				.LSULoadAccessFaultM(LSULoadAccessFaultM),
				.LSUStoreAmoAccessFaultM(LSUStoreAmoAccessFaultM),
				.LoadAccessFaultM(LoadAccessFaultM),
				.StoreAmoAccessFaultM(StoreAmoAccessFaultM),
				.HPTWInstrAccessFaultF(HPTWInstrAccessFaultF),
				.LoadPageFaultM(LoadPageFaultM),
				.StoreAmoPageFaultM(StoreAmoPageFaultM),
				.LSULoadPageFaultM(LSULoadPageFaultM),
				.LSUStoreAmoPageFaultM(LSUStoreAmoPageFaultM),
				.HPTWInstrPageFaultF(HPTWInstrPageFaultF)
			);
		end
		else begin : genblk3
			assign PreLSURWM = MemRWM;
			assign IHAdrM = IEUAdrExtM;
			assign LSUFunct3M = Funct3M;
			assign LSUFunct7M = Funct7M;
			assign LSUAtomicM = AtomicM;
			assign IHWriteDataM = WriteDataZM;
			assign LoadAccessFaultM = LSULoadAccessFaultM;
			assign StoreAmoAccessFaultM = LSUStoreAmoAccessFaultM;
			assign LoadPageFaultM = LSULoadPageFaultM;
			assign StoreAmoPageFaultM = LSUStoreAmoPageFaultM;
			assign {HPTWStall, SelHPTW, PTE, PageType, DTLBWriteM, ITLBWriteF, HPTWFlushW} = 1'sb0;
			assign {HPTWInstrAccessFaultF, HPTWInstrPageFaultF} = 1'sb0;
		end
	endgenerate
	assign CommittedM = (SelHPTW | DCacheCommittedM) | BusCommittedM;
	assign GatedStallW = StallW & ~SelHPTW;
	assign DCacheBusStallM = DCacheStallM | LSUBusStallM;
	assign CacheBusHPWTStall = DCacheBusStallM | HPTWStall;
	assign LSUStallM = CacheBusHPWTStall | SpillStallM;
	generate
		if (P[4086] == 1) begin : dmmu
			wire DisableTranslation;
			wire WriteAccessM;
			wire DataUpdateDAM;
			assign DisableTranslation = SelHPTW | FlushDCacheM;
			assign WriteAccessM = PreLSURWM[0];
			mmu #(
				.P(P),
				.TLB_ENTRIES($signed(P[4017-:32])),
				.IMMU(0)
			) dmmu(
				.clk(clk),
				.reset(reset),
				.SATP_REGW(SATP_REGW),
				.STATUS_MXR(STATUS_MXR),
				.STATUS_SUM(STATUS_SUM),
				.STATUS_MPRV(STATUS_MPRV),
				.STATUS_MPP(STATUS_MPP),
				.ENVCFG_PBMTE(ENVCFG_PBMTE),
				.ENVCFG_ADUE(ENVCFG_ADUE),
				.PrivilegeModeW(PrivilegeModeW),
				.DisableTranslation(DisableTranslation),
				.VAdr(IHAdrM),
				.Size(LSUFunct3M[1:0]),
				.PTE(PTE),
				.PageTypeWriteVal(PageType),
				.TLBWrite(DTLBWriteM),
				.TLBFlush(sfencevmaM),
				.PhysicalAddress(PAdrM),
				.TLBMiss(DTLBMissM),
				.Cacheable(CacheableM),
				.Idempotent(),
				.SelTIM(SelDTIM),
				.InstrAccessFaultF(),
				.LoadAccessFaultM(LSULoadAccessFaultM),
				.StoreAmoAccessFaultM(LSUStoreAmoAccessFaultM),
				.InstrPageFaultF(),
				.LoadPageFaultM(LSULoadPageFaultM),
				.StoreAmoPageFaultM(LSUStoreAmoPageFaultM),
				.LoadMisalignedFaultM(LoadMisalignedFaultM),
				.StoreAmoMisalignedFaultM(StoreAmoMisalignedFaultM),
				.UpdateDA(DataUpdateDAM),
				.CMOpM(CMOpM),
				.AtomicAccessM(|LSUAtomicM),
				.ExecuteAccessF(1'b0),
				.WriteAccessM(WriteAccessM),
				.ReadAccessM(PreLSURWM[1]),
				.PMPCFG_ARRAY_REGW(PMPCFG_ARRAY_REGW),
				.PMPADDR_ARRAY_REGW(PMPADDR_ARRAY_REGW)
			);
			assign DTLBMissOrUpdateDAM = DTLBMissM | (P[4064] & DataUpdateDAM);
		end
		else begin : genblk4
			assign DTLBMissOrUpdateDAM = 1'sb0;
			assign {DTLBMissM, LSULoadAccessFaultM, LSUStoreAmoAccessFaultM, LoadMisalignedFaultM, StoreAmoMisalignedFaultM} = 1'sb0;
			assign {LSULoadPageFaultM, LSUStoreAmoPageFaultM} = 1'sb0;
			assign PAdrM = IHAdrM[$signed(P[1640-:32]) - 1:0];
			assign CacheableM = 1'b1;
			assign SelDTIM = P[3600] & ~P[4052];
		end
	endgenerate
	assign LSUFlushW = HPTWFlushW | FlushW;
	generate
		if (P[3600]) begin : dtim
			wire [$signed(P[1640-:32]) - 1:0] DTIMAdr;
			wire [1:0] DTIMMemRWM;
			mux2 #(.WIDTH($signed(P[1640-:32]))) DTIMAdrMux(
				.d0(IEUAdrExtE[$signed(P[1640-:32]) - 1:0]),
				.d1(IEUAdrExtM[$signed(P[1640-:32]) - 1:0]),
				.s(MemRWM[0]),
				.y(DTIMAdr)
			);
			assign DTIMMemRWM = (SelDTIM ? LSURWM : 0);
			dtim #(.P(P)) dtim(
				.clk(clk),
				.reset(reset),
				.ce(~GatedStallW),
				.MemRWM(DTIMMemRWM),
				.DTIMAdr(DTIMAdr),
				.FlushW(LSUFlushW),
				.WriteDataM(LSUWriteDataM),
				.ReadDataWordM(DTIMReadDataWordM[$signed(P[383-:32]) - 1:0]),
				.ByteMaskM(ByteMaskM)
			);
		end
		else begin : genblk5
			assign DTIMReadDataWordM = 1'sb0;
		end
		if (P[4052]) begin : bus
			if (P[4051]) begin : dcache
				localparam LLENWORDSPERLINE = $signed(P[3921-:32]) / $signed(P[383-:32]);
				localparam LLENLOGBWPL = $clog2(LLENWORDSPERLINE);
				localparam BEATSPERLINE = $signed(P[3921-:32]) / $signed(P[4151-:32]);
				localparam AHBWLOGBWPL = $clog2(BEATSPERLINE);
				localparam LINELEN = $signed(P[3921-:32]);
				localparam LLENPOVERAHBW = $signed(P[383-:32]) / $signed(P[4151-:32]);
				localparam CACHEWORDLEN = (P[4059] ? 2 * $signed(P[383-:32]) : $signed(P[383-:32]));
				wire [LINELEN - 1:0] FetchBuffer;
				wire [$signed(P[1640-:32]) - 1:0] DCacheBusAdr;
				wire [AHBWLOGBWPL - 1:0] BeatCount;
				wire DCacheBusAck;
				wire SelBusBeat;
				wire [1:0] CacheBusRW;
				wire [1:0] BusRW;
				wire CacheableOrFlushCacheM;
				wire [1:0] CacheRWM;
				wire FlushDCache;
				wire BusCMOZero;
				wire [3:0] CacheCMOpM;
				wire BusAtomic;
				if (P[4061]) begin : genblk1
					assign BusCMOZero = CMOpM[3] & ~CacheableM;
					assign CacheCMOpM = (CacheableM & ~SelHPTW ? CMOpM : {4 {1'sb0}});
					assign BusAtomic = AtomicM[1] & ~CacheableM;
				end
				else begin : genblk1
					assign BusCMOZero = 1'b0;
					assign CacheCMOpM = 1'sb0;
					assign BusAtomic = 1'b0;
				end
				assign BusRW = (~CacheableM & ~SelDTIM ? LSURWM : {2 {1'sb0}});
				assign CacheableOrFlushCacheM = CacheableM | FlushDCacheM;
				assign CacheRWM = (CacheableM & ~SelDTIM ? LSURWM : {2 {1'sb0}});
				assign FlushDCache = FlushDCacheM & ~SelHPTW;
				cache #(
					.P(P),
					.PA_BITS($signed(P[1640-:32])),
					.LINELEN($signed(P[3921-:32])),
					.NUMSETS(($signed(P[3953-:32]) * 8) / LINELEN),
					.NUMWAYS($signed(P[3985-:32])),
					.LOGBWPL(LLENLOGBWPL),
					.WORDLEN(CACHEWORDLEN),
					.MUXINTERVAL($signed(P[383-:32])),
					.READ_ONLY_CACHE(0)
				) dcache(
					.clk(clk),
					.reset(reset),
					.Stall(GatedStallW & ~SelSpillE),
					.SelBusBeat(SelBusBeat),
					.FlushStage(LSUFlushW),
					.CacheRW(CacheRWM),
					.FlushCache(FlushDCache),
					.NextSet(IEUAdrExtE[11:0]),
					.PAdr(PAdrM),
					.ByteMask(ByteMaskSpillM),
					.BeatCount(BeatCount[AHBWLOGBWPL - 1:AHBWLOGBWPL - LLENLOGBWPL]),
					.WriteData(LSUWriteDataSpillM),
					.SelHPTW(SelHPTW),
					.CacheStall(DCacheStallM),
					.CacheMiss(DCacheMiss),
					.CacheAccess(DCacheAccess),
					.CacheCommitted(DCacheCommittedM),
					.CacheBusAdr(DCacheBusAdr),
					.ReadDataWord(DCacheReadDataWordM),
					.FetchBuffer(FetchBuffer),
					.CacheBusRW(CacheBusRW),
					.CacheBusAck(DCacheBusAck),
					.InvalidateCache(1'b0),
					.CMOpM(CacheCMOpM)
				);
				ahbcacheinterface #(
					.P(P),
					.BEATSPERLINE(BEATSPERLINE),
					.AHBWLOGBWPL(AHBWLOGBWPL),
					.LINELEN(LINELEN),
					.LLENPOVERAHBW(LLENPOVERAHBW),
					.READ_ONLY_CACHE(0)
				) ahbcacheinterface(
					.HCLK(clk),
					.HRESETn(~reset),
					.Flush(LSUFlushW),
					.HRDATA(HRDATA),
					.HWDATA(LSUHWDATA),
					.HWSTRB(LSUHWSTRB),
					.HSIZE(LSUHSIZE),
					.HBURST(LSUHBURST),
					.HTRANS(LSUHTRANS),
					.HWRITE(LSUHWRITE),
					.HREADY(LSUHREADY),
					.BeatCount(BeatCount),
					.SelBusBeat(SelBusBeat),
					.CacheReadDataWordM(DCacheReadDataWordM[$signed(P[383-:32]) - 1:0]),
					.WriteDataM(LSUWriteDataM),
					.Funct3(LSUFunct3M),
					.HADDR(LSUHADDR),
					.CacheBusAdr(DCacheBusAdr),
					.CacheBusRW(CacheBusRW),
					.BusAtomic(BusAtomic),
					.BusCMOZero(BusCMOZero),
					.CacheableOrFlushCacheM(CacheableOrFlushCacheM),
					.CacheBusAck(DCacheBusAck),
					.FetchBuffer(FetchBuffer),
					.PAdr(PAdrM),
					.Cacheable(CacheableOrFlushCacheM),
					.BusRW(BusRW),
					.Stall(GatedStallW),
					.BusStall(LSUBusStallM),
					.BusCommitted(BusCommittedM)
				);
				mux3 #(.WIDTH($signed(P[383-:32]))) UnCachedDataMux(
					.d0(DCacheReadDataWordSpillM),
					.d1({LLENPOVERAHBW {FetchBuffer[$signed(P[4216-:32]) - 1:0]}}),
					.d2({{$signed(P[383-:32]) - $signed(P[4216-:32]) {1'b0}}, DTIMReadDataWordM[$signed(P[4216-:32]) - 1:0]}),
					.s({SelDTIM, ~CacheableOrFlushCacheM}),
					.y(ReadDataWordMuxM)
				);
			end
			else begin : passthrough
				wire [1:0] BusRW;
				wire [$signed(P[4216-:32]) - 1:0] FetchBuffer;
				assign BusRW = (~SelDTIM ? LSURWM : 0);
				assign LSUHADDR = PAdrM;
				assign LSUHSIZE = LSUFunct3M;
				ahbinterface #(
					.XLEN($signed(P[4216-:32])),
					.LSU(1'b1)
				) ahbinterface(
					.HCLK(clk),
					.HRESETn(~reset),
					.Flush(LSUFlushW),
					.HREADY(LSUHREADY),
					.HRDATA(HRDATA),
					.HTRANS(LSUHTRANS),
					.HWRITE(LSUHWRITE),
					.HWDATA(LSUHWDATA),
					.HWSTRB(LSUHWSTRB),
					.BusRW(BusRW),
					.BusAtomic(AtomicM[1]),
					.ByteMask(ByteMaskM[($signed(P[4216-:32]) / 8) - 1:0]),
					.WriteData(LSUWriteDataM[$signed(P[4216-:32]) - 1:0]),
					.Stall(GatedStallW),
					.BusStall(LSUBusStallM),
					.BusCommitted(BusCommittedM),
					.FetchBuffer(FetchBuffer)
				);
				if (P[3600]) begin : genblk1
					mux2 #(.WIDTH($signed(P[4216-:32]))) ReadDataMux2(
						.d0(FetchBuffer),
						.d1(DTIMReadDataWordM[$signed(P[4216-:32]) - 1:0]),
						.s(SelDTIM),
						.y(ReadDataWordMuxM[$signed(P[4216-:32]) - 1:0])
					);
				end
				else begin : genblk1
					assign ReadDataWordMuxM[$signed(P[4216-:32]) - 1:0] = FetchBuffer[$signed(P[4216-:32]) - 1:0];
				end
				assign LSUHBURST = 3'b000;
				assign {DCacheStallM, DCacheCommittedM, DCacheMiss, DCacheAccess, DCacheReadDataWordM} = 1'sb0;
			end
		end
		else begin : nobus
			assign {LSUHWDATA, LSUHADDR, LSUHWRITE, LSUHSIZE, LSUHBURST, LSUHTRANS, LSUHWSTRB} = 1'sb0;
			assign DCacheReadDataWordM = 1'sb0;
			assign ReadDataWordMuxM = DTIMReadDataWordM;
			assign {LSUBusStallM, BusCommittedM} = 1'sb0;
			assign {DCacheMiss, DCacheAccess} = 1'sb0;
			assign {DCacheStallM, DCacheCommittedM} = 1'sb0;
		end
		if (P[4054] | P[4053]) begin : atomic
			atomic #(.P(P)) atomic(
				.clk(clk),
				.reset(reset),
				.StallW(StallW),
				.ReadDataM(ReadDataM[$signed(P[4216-:32]) - 1:0]),
				.IHWriteDataM(IHWriteDataM),
				.PAdrM(PAdrM),
				.LSUFunct7M(LSUFunct7M),
				.LSUFunct3M(LSUFunct3M),
				.LSUAtomicM(LSUAtomicM),
				.PreLSURWM(PreLSURWM),
				.LSUFlushW(LSUFlushW),
				.IMAWriteDataM(IMAWriteDataM),
				.SquashSCW(SquashSCW),
				.LSURWM(LSURWM)
			);
		end
		else begin : lrsc
			assign SquashSCW = 1'b0;
			assign LSURWM = PreLSURWM;
			assign IMAWriteDataM = IHWriteDataM;
		end
		if (P[1491]) begin : genblk8
			if ($signed(P[901-:32]) >= $signed(P[4216-:32])) begin : genblk1
				mux2 #(.WIDTH($signed(P[383-:32]))) datamux(
					.d0({{{$signed(P[383-:32]) - $signed(P[4216-:32])} {1'b0}}, IMAWriteDataM}),
					.d1(FWriteDataM),
					.s(FpLoadStoreM),
					.y(IMAFWriteDataM)
				);
			end
			else begin : genblk1
				mux2 #(.WIDTH($signed(P[383-:32]))) datamux(
					.d0(IMAWriteDataM),
					.d1({{{$signed(P[4216-:32]) - $signed(P[901-:32])} {1'b0}}, FWriteDataM}),
					.s(FpLoadStoreM),
					.y(IMAFWriteDataM)
				);
			end
		end
		else begin : genblk8
			assign IMAFWriteDataM = IMAWriteDataM;
		end
	endgenerate
	subwordread #(.P(P)) subwordread(
		.ReadDataWordMuxM(LittleEndianReadDataWordM),
		.PAdrM(PAdrM[3:0]),
		.BigEndianM(BigEndianM),
		.FpLoadStoreM(FpLoadStoreM),
		.Funct3M(LSUFunct3M),
		.ReadDataM(ReadDataM)
	);
	subwordwrite #(.LLEN($signed(P[383-:32]))) subwordwrite(
		.LSUFunct3M(LSUFunct3M),
		.IMAFWriteDataM(IMAFWriteDataM),
		.LittleEndianWriteDataM(LittleEndianWriteDataM)
	);
	swbytemask #(
		.WORDLEN($signed(P[383-:32])),
		.EXTEND(P[4059])
	) swbytemask(
		.Size(LSUFunct3M),
		.Adr(PAdrM[$clog2($signed(P[383-:32]) / 8) - 1:0]),
		.ByteMask(ByteMaskM),
		.ByteMaskExtended(ByteMaskExtendedM)
	);
	flopen #(.WIDTH($signed(P[383-:32]))) ReadDataMWReg(
		.clk(clk),
		.en(~StallW),
		.d(ReadDataM),
		.q(ReadDataW)
	);
	generate
		if (P[4065]) begin : endian
			endianswap #(.LEN($signed(P[383-:32]))) storeswap(
				.BigEndianM(BigEndianM),
				.a(LittleEndianWriteDataM),
				.y(LSUWriteDataM)
			);
			endianswap #(.LEN($signed(P[383-:32]))) loadswap(
				.BigEndianM(BigEndianM),
				.a(ReadDataWordMuxM),
				.y(LittleEndianReadDataWordM)
			);
		end
		else begin : genblk9
			assign LSUWriteDataM = LittleEndianWriteDataM;
			assign LittleEndianReadDataWordM = ReadDataWordMuxM;
		end
	endgenerate
endmodule
module subwordread (
	ReadDataWordMuxM,
	PAdrM,
	Funct3M,
	FpLoadStoreM,
	BigEndianM,
	ReadDataM
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[383-:32]) - 1:0] ReadDataWordMuxM;
	input wire [3:0] PAdrM;
	input wire [2:0] Funct3M;
	input wire FpLoadStoreM;
	input wire BigEndianM;
	output reg [$signed(P[383-:32]) - 1:0] ReadDataM;
	localparam ADRBITS = $clog2($signed(P[383-:32])) - 3;
	wire [ADRBITS - 1:0] PAdrSwapM;
	wire [7:0] ByteM;
	wire [15:0] HalfwordM;
	wire [31:0] WordM;
	wire [63:0] DblWordM;
	generate
		if (P[4065]) begin : genblk1
			assign PAdrSwapM = PAdrM[ADRBITS - 1:0] ^ {ADRBITS {BigEndianM}};
		end
		else begin : genblk1
			assign PAdrSwapM = PAdrM[ADRBITS - 1:0];
		end
		if ($signed(P[383-:32]) == 128) begin : genblk2
			mux2 #(.WIDTH(64)) dblmux(
				.d0(ReadDataWordMuxM[63:0]),
				.d1(ReadDataWordMuxM[127:64]),
				.s(PAdrSwapM[3]),
				.y(DblWordM)
			);
		end
		else if ($signed(P[383-:32]) == 64) begin : genblk2
			assign DblWordM = ReadDataWordMuxM;
		end
		else begin : genblk2
			assign DblWordM = 1'sb0;
		end
		if ($signed(P[383-:32]) >= 64) begin : genblk3
			mux2 #(.WIDTH(32)) wordmux(
				.d0(DblWordM[31:0]),
				.d1(DblWordM[63:32]),
				.s(PAdrSwapM[2]),
				.y(WordM)
			);
		end
		else begin : genblk3
			assign WordM = ReadDataWordMuxM;
		end
	endgenerate
	mux2 #(.WIDTH(16)) halfwordmux(
		.d0(WordM[15:0]),
		.d1(WordM[31:16]),
		.s(PAdrSwapM[1]),
		.y(HalfwordM)
	);
	mux2 #(.WIDTH(8)) bytemux(
		.d0(HalfwordM[7:0]),
		.d1(HalfwordM[15:8]),
		.s(PAdrSwapM[0]),
		.y(ByteM)
	);
	always @(*) begin
		if (_sv2v_0)
			;
		case (Funct3M)
			3'b000: ReadDataM = {{$signed(P[383-:32]) - 8 {ByteM[7]}}, ByteM};
			3'b001: ReadDataM = {{$signed(P[383-:32]) - 16 {HalfwordM[15] | FpLoadStoreM}}, HalfwordM[15:0]};
			3'b010: ReadDataM = {{$signed(P[383-:32]) - 32 {WordM[31] | FpLoadStoreM}}, WordM[31:0]};
			3'b011:
				if ($signed(P[383-:32]) >= 64)
					ReadDataM = {{$signed(P[383-:32]) - 64 {DblWordM[63] | FpLoadStoreM}}, DblWordM[63:0]};
				else
					ReadDataM = ReadDataWordMuxM;
			3'b100:
				if ($signed(P[383-:32]) == 128)
					ReadDataM = (FpLoadStoreM ? ReadDataWordMuxM : {{$signed(P[383-:32]) - 8 {1'b0}}, ByteM[7:0]});
				else
					ReadDataM = {{$signed(P[383-:32]) - 8 {1'b0}}, ByteM[7:0]};
			3'b101: ReadDataM = {{$signed(P[383-:32]) - 16 {1'b0}}, HalfwordM[15:0]};
			3'b110: ReadDataM = {{$signed(P[383-:32]) - 32 {1'b0}}, WordM[31:0]};
			default: ReadDataM = ReadDataWordMuxM;
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
module subwordwrite (
	LSUFunct3M,
	IMAFWriteDataM,
	LittleEndianWriteDataM
);
	reg _sv2v_0;
	parameter LLEN = 0;
	input wire [2:0] LSUFunct3M;
	input wire [LLEN - 1:0] IMAFWriteDataM;
	output reg [LLEN - 1:0] LittleEndianWriteDataM;
	generate
		if (LLEN == 128) begin : sww
			always @(*) begin
				if (_sv2v_0)
					;
				case (LSUFunct3M[2:0])
					3'b000: LittleEndianWriteDataM = {16 {IMAFWriteDataM[7:0]}};
					3'b001: LittleEndianWriteDataM = {8 {IMAFWriteDataM[15:0]}};
					3'b010: LittleEndianWriteDataM = {4 {IMAFWriteDataM[31:0]}};
					3'b011: LittleEndianWriteDataM = {2 {IMAFWriteDataM[63:0]}};
					default: LittleEndianWriteDataM = IMAFWriteDataM;
				endcase
			end
		end
		else if (LLEN == 64) begin : sww
			always @(*) begin
				if (_sv2v_0)
					;
				case (LSUFunct3M[1:0])
					2'b00: LittleEndianWriteDataM = {8 {IMAFWriteDataM[7:0]}};
					2'b01: LittleEndianWriteDataM = {4 {IMAFWriteDataM[15:0]}};
					2'b10: LittleEndianWriteDataM = {2 {IMAFWriteDataM[31:0]}};
					2'b11: LittleEndianWriteDataM = IMAFWriteDataM;
				endcase
			end
		end
		else begin : sww
			always @(*) begin
				if (_sv2v_0)
					;
				case (LSUFunct3M[1:0])
					2'b00: LittleEndianWriteDataM = {4 {IMAFWriteDataM[7:0]}};
					2'b01: LittleEndianWriteDataM = {2 {IMAFWriteDataM[15:0]}};
					2'b10: LittleEndianWriteDataM = IMAFWriteDataM;
					default: LittleEndianWriteDataM = IMAFWriteDataM;
				endcase
			end
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module swbytemask (
	Size,
	Adr,
	ByteMask,
	ByteMaskExtended
);
	parameter WORDLEN = 0;
	parameter EXTEND = 0;
	input wire [2:0] Size;
	input wire [$clog2(WORDLEN / 8) - 1:0] Adr;
	output wire [(WORDLEN / 8) - 1:0] ByteMask;
	output wire [(WORDLEN / 8) - 1:0] ByteMaskExtended;
	generate
		if (EXTEND) begin : genblk1
			wire [((WORDLEN * 2) / 8) - 1:0] ExtendedByteMask;
			assign ExtendedByteMask = (('d2 ** ('d2 ** Size)) - 'd1) << Adr;
			assign ByteMask = ExtendedByteMask[(WORDLEN / 8) - 1:0];
			assign ByteMaskExtended = ExtendedByteMask[((WORDLEN * 2) / 8) - 1:WORDLEN / 8];
		end
		else begin : genblk1
			assign ByteMask = (('d2 ** ('d2 ** Size)) - 'd1) << Adr;
			assign ByteMaskExtended = 1'sb0;
		end
	endgenerate
endmodule
module div (
	clk,
	reset,
	StallM,
	FlushE,
	IntDivE,
	DivSignedE,
	W64E,
	ForwardedSrcAE,
	ForwardedSrcBE,
	DivBusyE,
	QuotM,
	RemM
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallM;
	input wire FlushE;
	input wire IntDivE;
	input wire DivSignedE;
	input wire W64E;
	input wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcAE;
	input wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcBE;
	output wire DivBusyE;
	output wire [$signed(P[4216-:32]) - 1:0] QuotM;
	output wire [$signed(P[4216-:32]) - 1:0] RemM;
	localparam STEPBITS = $clog2($signed(P[4216-:32]) / $signed(P[3761-:32]));
	reg [1:0] state;
	wire [$signed(P[4216-:32]) - 1:0] W [$signed(P[3761-:32]):0];
	wire [$signed(P[4216-:32]) - 1:0] XQ [$signed(P[3761-:32]):0];
	wire [$signed(P[4216-:32]) - 1:0] WNext;
	wire [$signed(P[4216-:32]) - 1:0] XQNext;
	wire [$signed(P[4216-:32]) - 1:0] DinE;
	wire [$signed(P[4216-:32]) - 1:0] XinE;
	wire [$signed(P[4216-:32]) - 1:0] DnE;
	wire [$signed(P[4216-:32]) - 1:0] DAbsBE;
	wire [$signed(P[4216-:32]) - 1:0] DAbsB;
	wire [$signed(P[4216-:32]) - 1:0] XnE;
	wire [$signed(P[4216-:32]) - 1:0] XInitE;
	wire [$signed(P[4216-:32]) - 1:0] WnM;
	wire [$signed(P[4216-:32]) - 1:0] XQnM;
	reg [STEPBITS:0] step;
	wire Div0E;
	wire Div0M;
	wire DivStartE;
	wire SignXE;
	wire SignDE;
	wire NegQE;
	wire NegWM;
	wire NegQM;
	assign DivStartE = (IntDivE & (state == 2'd0)) & ~StallM;
	assign DivBusyE = (state == 2'd1) | DivStartE;
	generate
		if ($signed(P[4216-:32]) == 64) begin : rv64
			mux2 #(.WIDTH($signed(P[4216-:32]))) xinmux(
				.d0(ForwardedSrcAE),
				.d1({ForwardedSrcAE[31:0], 32'b00000000000000000000000000000000}),
				.s(W64E),
				.y(XinE)
			);
			mux2 #(.WIDTH($signed(P[4216-:32]))) dinmux(
				.d0(ForwardedSrcBE),
				.d1({{32 {ForwardedSrcBE[31] & DivSignedE}}, ForwardedSrcBE[31:0]}),
				.s(W64E),
				.y(DinE)
			);
		end
		else begin : genblk1
			assign XinE = ForwardedSrcAE;
			assign DinE = ForwardedSrcBE;
		end
	endgenerate
	assign SignDE = DivSignedE & DinE[$signed(P[4216-:32]) - 1];
	assign SignXE = DivSignedE & XinE[$signed(P[4216-:32]) - 1];
	assign NegQE = SignDE ^ SignXE;
	assign Div0E = DinE == 0;
	neg #(.WIDTH($signed(P[4216-:32]))) negd(
		.a(DinE),
		.y(DnE)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) dabsmux(
		.d0(DnE),
		.d1(DinE),
		.s(SignDE),
		.y(DAbsBE)
	);
	neg #(.WIDTH($signed(P[4216-:32]))) negx(
		.a(XinE),
		.y(XnE)
	);
	mux3 #(.WIDTH($signed(P[4216-:32]))) xabsmux(
		.d0(XinE),
		.d1(XnE),
		.d2(ForwardedSrcAE),
		.s({Div0E, SignXE}),
		.y(XInitE)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) wmux(
		.d0(W[$signed(P[3761-:32])]),
		.d1({$signed(P[4216-:32]) {1'b0}}),
		.s(DivStartE),
		.y(WNext)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) xmux(
		.d0(XQ[$signed(P[3761-:32])]),
		.d1(XInitE),
		.s(DivStartE),
		.y(XQNext)
	);
	flopen #(.WIDTH($signed(P[4216-:32]))) wreg(
		.clk(clk),
		.en(DivBusyE),
		.d(WNext),
		.q(W[0])
	);
	flopen #(.WIDTH($signed(P[4216-:32]))) xreg(
		.clk(clk),
		.en(DivBusyE),
		.d(XQNext),
		.q(XQ[0])
	);
	flopen #(.WIDTH($signed(P[4216-:32]))) dabsreg(
		.clk(clk),
		.en(DivStartE),
		.d(DAbsBE),
		.q(DAbsB)
	);
	genvar _gv_i_3;
	generate
		for (_gv_i_3 = 0; _gv_i_3 < $signed(P[3761-:32]); _gv_i_3 = _gv_i_3 + 1) begin : genblk2
			localparam i = _gv_i_3;
			divstep #(.XLEN($signed(P[4216-:32]))) divstep(
				.W(W[i]),
				.XQ(XQ[i]),
				.DAbsB(DAbsB),
				.WOut(W[i + 1]),
				.XQOut(XQ[i + 1])
			);
		end
	endgenerate
	flopen #(.WIDTH(3)) Div0eMReg(
		.clk(clk),
		.en(DivStartE),
		.d({Div0E, NegQE, SignXE}),
		.q({Div0M, NegQM, NegWM})
	);
	neg #(.WIDTH($signed(P[4216-:32]))) qneg(
		.a(XQ[0]),
		.y(XQnM)
	);
	neg #(.WIDTH($signed(P[4216-:32]))) wneg(
		.a(W[0]),
		.y(WnM)
	);
	mux3 #(.WIDTH($signed(P[4216-:32]))) qmux(
		.d0(XQ[0]),
		.d1(XQnM),
		.d2({$signed(P[4216-:32]) {1'b1}}),
		.s({Div0M, NegQM}),
		.y(QuotM)
	);
	mux3 #(.WIDTH($signed(P[4216-:32]))) remmux(
		.d0(W[0]),
		.d1(WnM),
		.d2(XQ[0]),
		.s({Div0M, NegWM}),
		.y(RemM)
	);
	always @(posedge clk)
		if (reset | FlushE)
			state <= 2'd0;
		else if (DivStartE) begin
			step <= 1;
			if (Div0E)
				state <= 2'd2;
			else
				state <= 2'd1;
		end
		else if (state == 2'd1) begin
			if (step[STEPBITS] | ((($signed(P[4216-:32]) == 64) & W64E) & step[STEPBITS - 1]))
				state <= 2'd2;
			step <= step + 1;
		end
		else if (state == 2'd2) begin
			if (StallM)
				state <= 2'd2;
			else
				state <= 2'd0;
		end
endmodule
module divstep (
	W,
	XQ,
	DAbsB,
	WOut,
	XQOut
);
	parameter XLEN = 0;
	input wire [XLEN - 1:0] W;
	input wire [XLEN - 1:0] XQ;
	input wire [XLEN - 1:0] DAbsB;
	output wire [XLEN - 1:0] WOut;
	output wire [XLEN - 1:0] XQOut;
	wire [XLEN - 1:0] WShift;
	wire [XLEN - 1:0] WPrime;
	wire qi;
	wire qib;
	assign {WShift, XQOut} = {W[XLEN - 2:0], XQ, qi};
	adder #(.WIDTH(XLEN + 1)) wdsub(
		.a({1'b0, WShift}),
		.b({1'b1, DAbsB}),
		.y({qib, WPrime})
	);
	assign qi = ~qib;
	mux2 #(.WIDTH(XLEN)) wrestoremux(
		.d0(WShift),
		.d1(WPrime),
		.s(qi),
		.y(WOut)
	);
endmodule
module mdu (
	clk,
	reset,
	StallM,
	StallW,
	FlushE,
	FlushM,
	FlushW,
	ForwardedSrcAE,
	ForwardedSrcBE,
	Funct3E,
	Funct3M,
	IntDivE,
	W64E,
	MDUActiveE,
	MDUResultW,
	DivBusyE
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallM;
	input wire StallW;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	input wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcAE;
	input wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcBE;
	input wire [2:0] Funct3E;
	input wire [2:0] Funct3M;
	input wire IntDivE;
	input wire W64E;
	input wire MDUActiveE;
	output wire [$signed(P[4216-:32]) - 1:0] MDUResultW;
	output wire DivBusyE;
	wire [($signed(P[4216-:32]) * 2) - 1:0] ProdM;
	wire [$signed(P[4216-:32]) - 1:0] QuotM;
	wire [$signed(P[4216-:32]) - 1:0] RemM;
	reg [$signed(P[4216-:32]) - 1:0] PrelimResultM;
	wire [$signed(P[4216-:32]) - 1:0] MDUResultM;
	wire W64M;
	mul #(.XLEN($signed(P[4216-:32]))) mul(
		.clk(clk),
		.reset(reset),
		.StallM(StallM),
		.FlushM(FlushM),
		.ForwardedSrcAE(ForwardedSrcAE),
		.ForwardedSrcBE(ForwardedSrcBE),
		.Funct3E(Funct3E),
		.ProdM(ProdM)
	);
	generate
		if ((P[3729] & P[1491]) | !P[1489]) begin : nodiv
			assign QuotM = 1'sb0;
			assign RemM = 1'sb0;
			assign DivBusyE = 1'b0;
		end
		else begin : div
			div #(.P(P)) div(
				.clk(clk),
				.reset(reset),
				.StallM(StallM),
				.FlushE(FlushE),
				.DivSignedE(~Funct3E[0]),
				.W64E(W64E),
				.IntDivE(IntDivE),
				.ForwardedSrcAE(ForwardedSrcAE),
				.ForwardedSrcBE(ForwardedSrcBE),
				.DivBusyE(DivBusyE),
				.QuotM(QuotM),
				.RemM(RemM)
			);
		end
	endgenerate
	always @(*) begin
		if (_sv2v_0)
			;
		case (Funct3M)
			3'b000: PrelimResultM = ProdM[$signed(P[4216-:32]) - 1:0];
			3'b001: PrelimResultM = ProdM[($signed(P[4216-:32]) * 2) - 1:$signed(P[4216-:32])];
			3'b010: PrelimResultM = ProdM[($signed(P[4216-:32]) * 2) - 1:$signed(P[4216-:32])];
			3'b011: PrelimResultM = ProdM[($signed(P[4216-:32]) * 2) - 1:$signed(P[4216-:32])];
			3'b100: PrelimResultM = QuotM;
			3'b101: PrelimResultM = QuotM;
			3'b110: PrelimResultM = RemM;
			3'b111: PrelimResultM = RemM;
		endcase
	end
	flopenrc #(.WIDTH(1)) W64MReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(W64E),
		.q(W64M)
	);
	generate
		if ($signed(P[4216-:32]) == 64) begin : resmux
			assign MDUResultM = (W64M ? {{32 {PrelimResultM[31]}}, PrelimResultM[31:0]} : PrelimResultM);
		end
		else begin : resmux
			assign MDUResultM = PrelimResultM;
		end
	endgenerate
	flopenrc #(.WIDTH($signed(P[4216-:32]))) MDUResultWReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(MDUResultM),
		.q(MDUResultW)
	);
	initial _sv2v_0 = 0;
endmodule
module mul (
	clk,
	reset,
	StallM,
	FlushM,
	ForwardedSrcAE,
	ForwardedSrcBE,
	Funct3E,
	ProdM
);
	reg _sv2v_0;
	parameter XLEN = 0;
	input wire clk;
	input wire reset;
	input wire StallM;
	input wire FlushM;
	input wire [XLEN - 1:0] ForwardedSrcAE;
	input wire [XLEN - 1:0] ForwardedSrcBE;
	input wire [2:0] Funct3E;
	output wire [(XLEN * 2) - 1:0] ProdM;
	wire [XLEN - 1:0] Aprime;
	wire [XLEN - 1:0] Bprime;
	wire MULH;
	wire MULHSU;
	wire [XLEN - 2:0] PA;
	wire [XLEN - 2:0] PB;
	wire PP;
	wire [(XLEN * 2) - 1:0] PP1E;
	wire [(XLEN * 2) - 1:0] PP2E;
	wire [(XLEN * 2) - 1:0] PP3E;
	reg [(XLEN * 2) - 1:0] PP4E;
	wire [(XLEN * 2) - 1:0] PP1M;
	wire [(XLEN * 2) - 1:0] PP2M;
	wire [(XLEN * 2) - 1:0] PP3M;
	wire [(XLEN * 2) - 1:0] PP4M;
	assign Aprime = {1'b0, ForwardedSrcAE[XLEN - 2:0]};
	assign Bprime = {1'b0, ForwardedSrcBE[XLEN - 2:0]};
	assign PP1E = Aprime * Bprime;
	assign PA = {XLEN - 1 {ForwardedSrcAE[XLEN - 1]}} & ForwardedSrcBE[XLEN - 2:0];
	assign PB = {XLEN - 1 {ForwardedSrcBE[XLEN - 1]}} & ForwardedSrcAE[XLEN - 2:0];
	assign PP = ForwardedSrcAE[XLEN - 1] & ForwardedSrcBE[XLEN - 1];
	assign MULH = Funct3E == 3'b001;
	assign MULHSU = Funct3E == 3'b010;
	assign PP2E = {2'b00, (MULH | MULHSU ? ~PA : PA), {XLEN - 1 {1'b0}}};
	assign PP3E = {2'b00, (MULH ? ~PB : PB), {XLEN - 1 {1'b0}}};
	always @(*) begin
		if (_sv2v_0)
			;
		if (MULH)
			PP4E = {1'b1, PP, {XLEN - 3 {1'b0}}, 1'b1, {XLEN {1'b0}}};
		else if (MULHSU)
			PP4E = {1'b1, ~PP, {XLEN - 2 {1'b0}}, 1'b1, {XLEN - 1 {1'b0}}};
		else
			PP4E = {1'b0, PP, {(XLEN * 2) - 2 {1'b0}}};
	end
	flopenrc #(.WIDTH(XLEN * 2)) PP1Reg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(PP1E),
		.q(PP1M)
	);
	flopenrc #(.WIDTH(XLEN * 2)) PP2Reg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(PP2E),
		.q(PP2M)
	);
	flopenrc #(.WIDTH(XLEN * 2)) PP3Reg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(PP3E),
		.q(PP3M)
	);
	flopenrc #(.WIDTH(XLEN * 2)) PP4Reg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(PP4E),
		.q(PP4M)
	);
	assign ProdM = ((PP1M + PP2M) + PP3M) + PP4M;
	initial _sv2v_0 = 0;
endmodule
module adrdec (
	PhysicalAddress,
	Base,
	Range,
	Supported,
	AccessValid,
	Size,
	SizeMask,
	Sel
);
	parameter PA_BITS = 0;
	input wire [PA_BITS - 1:0] PhysicalAddress;
	input wire [PA_BITS - 1:0] Base;
	input wire [PA_BITS - 1:0] Range;
	input wire Supported;
	input wire AccessValid;
	input wire [1:0] Size;
	input wire [3:0] SizeMask;
	output wire Sel;
	wire Match;
	wire SizeValid;
	assign Match = &((PhysicalAddress ~^ Base) | Range);
	assign SizeValid = SizeMask[Size];
	assign Sel = ((Match & Supported) & AccessValid) & SizeValid;
endmodule
module adrdecs (
	PhysicalAddress,
	AccessRW,
	AccessRX,
	AccessRWXC,
	Size,
	SelRegions
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[1640-:32]) - 1:0] PhysicalAddress;
	input wire AccessRW;
	input wire AccessRX;
	input wire AccessRWXC;
	input wire [1:0] Size;
	output wire [11:0] SelRegions;
	localparam [3:0] SUPPORTED_SIZE = ($signed(P[383-:32]) == 32 ? 4'b0111 : 4'b1111);
	adrdec #(.PA_BITS($signed(P[1640-:32]))) dtimdec(
		.PhysicalAddress(PhysicalAddress),
		.Base(P[3535 + $signed(P[1640-:32]):3536]),
		.Range(P[$signed(P[1640-:32]) + 3471:3472]),
		.Supported(P[3600]),
		.AccessValid(AccessRW),
		.Size(Size),
		.SizeMask(SUPPORTED_SIZE),
		.Sel(SelRegions[1])
	);
	adrdec #(.PA_BITS($signed(P[1640-:32]))) iromdec(
		.PhysicalAddress(PhysicalAddress),
		.Base(P[$signed(P[1640-:32]) + 3406:3407]),
		.Range(P[3342 + $signed(P[1640-:32]):3343]),
		.Supported(P[3471]),
		.AccessValid(AccessRX),
		.Size(Size),
		.SizeMask(SUPPORTED_SIZE),
		.Sel(SelRegions[2])
	);
	adrdec #(.PA_BITS($signed(P[1640-:32]))) ddr4dec(
		.PhysicalAddress(PhysicalAddress),
		.Base(P[3017 + $signed(P[1640-:32]):3018]),
		.Range(P[$signed(P[1640-:32]) + 2953:2954]),
		.Supported(P[3082]),
		.AccessValid(AccessRWXC),
		.Size(Size),
		.SizeMask(SUPPORTED_SIZE),
		.Sel(SelRegions[3])
	);
	adrdec #(.PA_BITS($signed(P[1640-:32]))) bootromdec(
		.PhysicalAddress(PhysicalAddress),
		.Base(P[3277 + $signed(P[1640-:32]):3278]),
		.Range(P[$signed(P[1640-:32]) + 3213:3214]),
		.Supported(P[3342]),
		.AccessValid(AccessRX),
		.Size(Size),
		.SizeMask(SUPPORTED_SIZE),
		.Sel(SelRegions[4])
	);
	adrdec #(.PA_BITS($signed(P[1640-:32]))) uncoreramdec(
		.PhysicalAddress(PhysicalAddress),
		.Base(P[3147 + $signed(P[1640-:32]):3148]),
		.Range(P[$signed(P[1640-:32]) + 3083:3084]),
		.Supported(P[3212]),
		.AccessValid(AccessRWXC),
		.Size(Size),
		.SizeMask(SUPPORTED_SIZE),
		.Sel(SelRegions[5])
	);
	adrdec #(.PA_BITS($signed(P[1640-:32]))) clintdec(
		.PhysicalAddress(PhysicalAddress),
		.Base(P[$signed(P[1640-:32]) + 2888:2889]),
		.Range(P[2824 + $signed(P[1640-:32]):2825]),
		.Supported(P[2953]),
		.AccessValid(AccessRW),
		.Size(Size),
		.SizeMask(SUPPORTED_SIZE),
		.Sel(SelRegions[6])
	);
	adrdec #(.PA_BITS($signed(P[1640-:32]))) gpiodec(
		.PhysicalAddress(PhysicalAddress),
		.Base(P[2759 + $signed(P[1640-:32]):2760]),
		.Range(P[$signed(P[1640-:32]) + 2695:2696]),
		.Supported(P[2824]),
		.AccessValid(AccessRW),
		.Size(Size),
		.SizeMask(4'b0100),
		.Sel(SelRegions[7])
	);
	adrdec #(.PA_BITS($signed(P[1640-:32]))) uartdec(
		.PhysicalAddress(PhysicalAddress),
		.Base(P[$signed(P[1640-:32]) + 2630:2631]),
		.Range(P[2566 + $signed(P[1640-:32]):2567]),
		.Supported(P[2695]),
		.AccessValid(AccessRW),
		.Size(Size),
		.SizeMask(4'b0001),
		.Sel(SelRegions[8])
	);
	adrdec #(.PA_BITS($signed(P[1640-:32]))) plicdec(
		.PhysicalAddress(PhysicalAddress),
		.Base(P[2501 + $signed(P[1640-:32]):2502]),
		.Range(P[$signed(P[1640-:32]) + 2437:2438]),
		.Supported(P[2566]),
		.AccessValid(AccessRW),
		.Size(Size),
		.SizeMask(4'b0100),
		.Sel(SelRegions[9])
	);
	adrdec #(.PA_BITS($signed(P[1640-:32]))) sdcdec(
		.PhysicalAddress(PhysicalAddress),
		.Base(P[$signed(P[1640-:32]) + 2372:2373]),
		.Range(P[2308 + $signed(P[1640-:32]):2309]),
		.Supported(P[2437]),
		.AccessValid(AccessRW),
		.Size(Size),
		.SizeMask(SUPPORTED_SIZE & 4'b1100),
		.Sel(SelRegions[10])
	);
	adrdec #(.PA_BITS($signed(P[1640-:32]))) spidec(
		.PhysicalAddress(PhysicalAddress),
		.Base(P[2243 + $signed(P[1640-:32]):2244]),
		.Range(P[$signed(P[1640-:32]) + 2179:2180]),
		.Supported(P[2308]),
		.AccessValid(AccessRW),
		.Size(Size),
		.SizeMask(4'b0100),
		.Sel(SelRegions[11])
	);
	assign SelRegions[0] = ~|SelRegions[11:1];
endmodule
module hptw (
	clk,
	reset,
	SATP_REGW,
	PCSpillF,
	IEUAdrExtM,
	MemRWM,
	AtomicM,
	STATUS_MXR,
	STATUS_SUM,
	STATUS_MPRV,
	STATUS_MPP,
	ENVCFG_ADUE,
	PrivilegeModeW,
	ReadDataM,
	WriteDataM,
	DCacheBusStallM,
	Funct3M,
	Funct7M,
	ITLBMissOrUpdateAF,
	DTLBMissOrUpdateDAM,
	FlushW,
	PTE,
	PageType,
	ITLBWriteF,
	DTLBWriteM,
	PreLSURWM,
	IHAdrM,
	IHWriteDataM,
	LSUAtomicM,
	LSUFunct3M,
	LSUFunct7M,
	HPTWFlushW,
	SelHPTW,
	HPTWStall,
	LSULoadAccessFaultM,
	LSUStoreAmoAccessFaultM,
	LSULoadPageFaultM,
	LSUStoreAmoPageFaultM,
	LoadAccessFaultM,
	StoreAmoAccessFaultM,
	HPTWInstrAccessFaultF,
	LoadPageFaultM,
	StoreAmoPageFaultM,
	HPTWInstrPageFaultF
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire [$signed(P[4216-:32]) - 1:0] SATP_REGW;
	input wire [$signed(P[4216-:32]) - 1:0] PCSpillF;
	input wire [$signed(P[4216-:32]) + 1:0] IEUAdrExtM;
	input wire [1:0] MemRWM;
	input wire [1:0] AtomicM;
	input wire STATUS_MXR;
	input wire STATUS_SUM;
	input wire STATUS_MPRV;
	input wire [1:0] STATUS_MPP;
	input wire ENVCFG_ADUE;
	input wire [1:0] PrivilegeModeW;
	input wire [$signed(P[4216-:32]) - 1:0] ReadDataM;
	input wire [$signed(P[4216-:32]) - 1:0] WriteDataM;
	input wire DCacheBusStallM;
	input wire [2:0] Funct3M;
	input wire [6:0] Funct7M;
	input wire ITLBMissOrUpdateAF;
	input wire DTLBMissOrUpdateDAM;
	input wire FlushW;
	output wire [$signed(P[4216-:32]) - 1:0] PTE;
	output wire [1:0] PageType;
	output wire ITLBWriteF;
	output wire DTLBWriteM;
	output wire [1:0] PreLSURWM;
	output wire [$signed(P[4216-:32]) + 1:0] IHAdrM;
	output wire [$signed(P[4216-:32]) - 1:0] IHWriteDataM;
	output wire [1:0] LSUAtomicM;
	output wire [2:0] LSUFunct3M;
	output wire [6:0] LSUFunct7M;
	output wire HPTWFlushW;
	output wire SelHPTW;
	output wire HPTWStall;
	input wire LSULoadAccessFaultM;
	input wire LSUStoreAmoAccessFaultM;
	input wire LSULoadPageFaultM;
	input wire LSUStoreAmoPageFaultM;
	output wire LoadAccessFaultM;
	output wire StoreAmoAccessFaultM;
	output wire HPTWInstrAccessFaultF;
	output wire LoadPageFaultM;
	output wire StoreAmoPageFaultM;
	output wire HPTWInstrPageFaultF;
	wire DTLBWalk;
	wire [$signed(P[1672-:32]) - 1:0] BasePageTablePPN;
	wire [$signed(P[1672-:32]) - 1:0] CurrentPPN;
	wire Executable;
	wire Writable;
	wire Readable;
	wire Valid;
	wire PTE_U;
	wire Misaligned;
	wire MegapageMisaligned;
	wire ValidPTE;
	wire LeafPTE;
	wire ValidLeafPTE;
	wire ValidNonLeafPTE;
	wire StartWalk;
	wire TLBMissOrUpdateDA;
	wire PRegEn;
	reg [1:0] NextPageType;
	wire [$signed(P[1608-:32]) - 1:0] SvMode;
	wire [$signed(P[4216-:32]) - 1:0] TranslationVAdr;
	wire [$signed(P[4216-:32]) - 1:0] NextPTE;
	wire [$signed(P[4216-:32]) - 1:0] NextPTE2;
	wire UpdatePTE;
	wire HPTWUpdateDA;
	wire [$signed(P[1640-:32]) - 1:0] HPTWReadAdr;
	wire SelHPTWAdr;
	wire [$signed(P[4216-:32]) + 1:0] HPTWAdrExt;
	wire LSUAccessFaultM;
	wire [$signed(P[1640-:32]) - 1:0] HPTWAdr;
	wire [1:0] HPTWRW;
	wire [2:0] HPTWSize;
	wire [3:0] WalkerState;
	reg [3:0] NextWalkerState;
	wire [3:0] InitialWalkerState;
	wire HPTWLoadAccessFault;
	wire HPTWStoreAmoAccessFault;
	wire HPTWInstrAccessFault;
	wire HPTWLoadAccessFaultDelay;
	wire HPTWStoreAmoAccessFaultDelay;
	wire HPTWInstrAccessFaultDelay;
	wire HPTWLoadPageFault;
	wire HPTWStoreAmoPageFault;
	wire HPTWInstrPageFault;
	wire HPTWLoadPageFaultDelay;
	wire HPTWStoreAmoPageFaultDelay;
	wire HPTWInstrPageFaultDelay;
	wire HPTWAccessFaultDelay;
	wire TakeHPTWFault;
	wire PBMTFaultM;
	wire DAUFaultM;
	wire PBMTOrDAUFaultM;
	wire HPTWFaultM;
	assign LSUAccessFaultM = LSULoadAccessFaultM | LSUStoreAmoAccessFaultM;
	assign PBMTOrDAUFaultM = PBMTFaultM | DAUFaultM;
	assign HPTWFaultM = LSUAccessFaultM | PBMTOrDAUFaultM;
	assign HPTWLoadAccessFault = ((LSUAccessFaultM & DTLBWalk) & MemRWM[1]) & ~MemRWM[0];
	assign HPTWStoreAmoAccessFault = (LSUAccessFaultM & DTLBWalk) & MemRWM[0];
	assign HPTWInstrAccessFault = LSUAccessFaultM & ~DTLBWalk;
	assign HPTWLoadPageFault = ((PBMTOrDAUFaultM & DTLBWalk) & MemRWM[1]) & ~MemRWM[0];
	assign HPTWStoreAmoPageFault = (PBMTOrDAUFaultM & DTLBWalk) & MemRWM[0];
	assign HPTWInstrPageFault = PBMTOrDAUFaultM & ~DTLBWalk;
	flopr #(.WIDTH(6)) HPTWAccesFaultReg(
		.clk(clk),
		.reset(reset),
		.d({HPTWLoadAccessFault, HPTWStoreAmoAccessFault, HPTWInstrAccessFault, HPTWLoadPageFault, HPTWStoreAmoPageFault, HPTWInstrPageFault}),
		.q({HPTWLoadAccessFaultDelay, HPTWStoreAmoAccessFaultDelay, HPTWInstrAccessFaultDelay, HPTWLoadPageFaultDelay, HPTWStoreAmoPageFaultDelay, HPTWInstrPageFaultDelay})
	);
	assign TakeHPTWFault = WalkerState != 4'd9;
	assign LoadAccessFaultM = (TakeHPTWFault ? HPTWLoadAccessFaultDelay : LSULoadAccessFaultM);
	assign StoreAmoAccessFaultM = (TakeHPTWFault ? HPTWStoreAmoAccessFaultDelay : LSUStoreAmoAccessFaultM);
	assign HPTWInstrAccessFaultF = (TakeHPTWFault ? HPTWInstrAccessFaultDelay : 1'b0);
	assign LoadPageFaultM = (TakeHPTWFault ? HPTWLoadPageFaultDelay : LSULoadPageFaultM);
	assign StoreAmoPageFaultM = (TakeHPTWFault ? HPTWStoreAmoPageFaultDelay : LSUStoreAmoPageFaultM);
	assign HPTWInstrPageFaultF = (TakeHPTWFault ? HPTWInstrPageFaultDelay : 1'b0);
	assign SvMode = SATP_REGW[$signed(P[4216-:32]) - 1:$signed(P[4216-:32]) - $signed(P[1608-:32])];
	assign BasePageTablePPN = SATP_REGW[$signed(P[1672-:32]) - 1:0];
	assign TLBMissOrUpdateDA = DTLBMissOrUpdateDAM | ITLBMissOrUpdateAF;
	mux2 #(.WIDTH($signed(P[4216-:32]))) vadrmux(
		.d0(PCSpillF),
		.d1(IEUAdrExtM[$signed(P[4216-:32]) - 1:0]),
		.s(DTLBWalk),
		.y(TranslationVAdr)
	);
	assign CurrentPPN = PTE[$signed(P[1672-:32]) + 9:10];
	flopenr #(.WIDTH(1)) TLBMissMReg(
		.clk(clk),
		.reset(reset),
		.en(StartWalk),
		.d(DTLBMissOrUpdateDAM),
		.q(DTLBWalk)
	);
	assign PRegEn = ((HPTWRW[1] & ~DCacheBusStallM) | UpdatePTE) | (NextWalkerState == 4'd9);
	assign NextPTE2 = (NextWalkerState == 4'd9 ? {$signed(P[4216-:32]) {1'sb0}} : NextPTE);
	flopenr #(.WIDTH($signed(P[4216-:32]))) PTEReg(
		.clk(clk),
		.reset(reset),
		.en(PRegEn),
		.d(NextPTE2),
		.q(PTE)
	);
	assign {PTE_U, Executable, Writable, Readable, Valid} = PTE[4:0];
	assign LeafPTE = (Executable | Writable) | Readable;
	assign ValidPTE = Valid & ~(Writable & ~Readable);
	assign ValidLeafPTE = ValidPTE & LeafPTE;
	assign ValidNonLeafPTE = Valid & ~LeafPTE;
	generate
		if ($signed(P[4216-:32]) == 64) begin : genblk1
			assign PBMTFaultM = ValidNonLeafPTE & |PTE[62:61];
		end
		else begin : genblk1
			assign PBMTFaultM = 1'b0;
		end
	endgenerate
	assign DAUFaultM = ValidNonLeafPTE & (|PTE[7:6] | PTE[4]);
	generate
		if (P[4064]) begin : hptwwrites
			wire ReadAccess;
			wire WriteAccess;
			wire InvalidRead;
			wire InvalidWrite;
			wire InvalidOp;
			wire UpperBitsUnequal;
			wire UpperBitsUnequalD;
			wire OtherPageFault;
			wire [1:0] EffectivePrivilegeMode;
			wire ImproperPrivilege;
			wire SaveHPTWAdr;
			wire SelHPTWWriteAdr;
			wire [$signed(P[1640-:32]) - 1:0] HPTWWriteAdr;
			wire SetDirty;
			wire Dirty;
			wire Accessed;
			wire [$signed(P[4216-:32]) - 1:0] AccessedPTE;
			assign AccessedPTE = {PTE[$signed(P[4216-:32]) - 1:8], SetDirty | PTE[7], 1'b1, PTE[5:0]};
			mux2 #(.WIDTH($signed(P[4216-:32]))) NextPTEMux(
				.d0(ReadDataM),
				.d1(AccessedPTE),
				.s(UpdatePTE),
				.y(NextPTE)
			);
			flopenr #(.WIDTH($signed(P[1640-:32]))) HPTWAdrWriteReg(
				.clk(clk),
				.reset(reset),
				.en(SaveHPTWAdr),
				.d(HPTWReadAdr),
				.q(HPTWWriteAdr)
			);
			assign SaveHPTWAdr = (((NextWalkerState == 4'd1) | (NextWalkerState == 4'd3)) | (NextWalkerState == 4'd5)) | (NextWalkerState == 4'd7);
			assign SelHPTWWriteAdr = UpdatePTE | HPTWRW[0];
			mux2 #(.WIDTH($signed(P[1640-:32]))) HPTWWriteAdrMux(
				.d0(HPTWReadAdr),
				.d1(HPTWWriteAdr),
				.s(SelHPTWWriteAdr),
				.y(HPTWAdr)
			);
			assign {Dirty, Accessed} = PTE[7:6];
			assign WriteAccess = MemRWM[0];
			assign SetDirty = (~Dirty & DTLBWalk) & WriteAccess;
			assign ReadAccess = MemRWM[1];
			assign EffectivePrivilegeMode = (DTLBWalk ? (STATUS_MPRV ? STATUS_MPP : PrivilegeModeW) : PrivilegeModeW);
			assign ImproperPrivilege = ((EffectivePrivilegeMode == P[1738-:2]) & ~PTE_U) | (((EffectivePrivilegeMode == P[1740-:2]) & PTE_U) & (~STATUS_SUM & DTLBWalk));
			vm64check #(.P(P)) vm64check(
				.SATP_MODE(SATP_REGW[$signed(P[4216-:32]) - 1:$signed(P[4216-:32]) - $signed(P[1608-:32])]),
				.VAdr(TranslationVAdr),
				.SV39Mode(),
				.UpperBitsUnequal(UpperBitsUnequal)
			);
			flopr #(.WIDTH(1)) upperbitsunequalreg(
				.clk(clk),
				.reset(reset),
				.d(UpperBitsUnequal),
				.q(UpperBitsUnequalD)
			);
			assign InvalidRead = (ReadAccess & ~Readable) & (~STATUS_MXR | ~Executable);
			assign InvalidWrite = WriteAccess & ~Writable;
			assign InvalidOp = (DTLBWalk ? InvalidRead | InvalidWrite : ~Executable);
			assign OtherPageFault = (((ImproperPrivilege | InvalidOp) | UpperBitsUnequalD) | Misaligned) | ~Valid;
			assign HPTWUpdateDA = ((ValidLeafPTE & (~Accessed | SetDirty)) & ENVCFG_ADUE) & ~OtherPageFault;
			assign HPTWRW[0] = WalkerState == 4'd10;
			assign UpdatePTE = (WalkerState == 4'd8) & HPTWUpdateDA;
		end
		else begin : genblk2
			assign NextPTE = ReadDataM;
			assign HPTWAdr = HPTWReadAdr;
			assign HPTWUpdateDA = 1'b0;
			assign UpdatePTE = 1'b0;
			assign HPTWRW[0] = 1'b0;
		end
	endgenerate
	assign StartWalk = (WalkerState == 4'd9) & TLBMissOrUpdateDA;
	assign HPTWRW[1] = (((WalkerState == 4'd7) | (WalkerState == 4'd5)) | (WalkerState == 4'd3)) | (WalkerState == 4'd1);
	assign DTLBWriteM = ((WalkerState == 4'd8) & ~HPTWUpdateDA) & DTLBWalk;
	assign ITLBWriteF = ((WalkerState == 4'd8) & ~HPTWUpdateDA) & ~DTLBWalk;
	flopr #(.WIDTH(2)) PageTypeReg(
		.clk(clk),
		.reset(reset),
		.d(NextPageType),
		.q(PageType)
	);
	always @(*) begin
		if (_sv2v_0)
			;
		case (WalkerState)
			4'd7: NextPageType = 2'b11;
			4'd5: NextPageType = 2'b10;
			4'd3: NextPageType = 2'b01;
			4'd1: NextPageType = 2'b00;
			default: NextPageType = PageType;
		endcase
	end
	generate
		if ($signed(P[4216-:32]) == 32) begin : genblk3
			reg [9:0] VPN;
			wire [$signed(P[1672-:32]) - 1:0] PPN;
			wire [10:1] sv2v_tmp_C200C;
			assign sv2v_tmp_C200C = ((WalkerState == 4'd2) | (WalkerState == 4'd3) ? TranslationVAdr[31:22] : TranslationVAdr[21:12]);
			always @(*) VPN = sv2v_tmp_C200C;
			assign PPN = ((WalkerState == 4'd2) | (WalkerState == 4'd3) ? BasePageTablePPN : CurrentPPN);
			assign HPTWReadAdr = {PPN, VPN, 2'b00};
			assign HPTWSize = 3'b010;
		end
		else begin : genblk3
			reg [8:0] VPN;
			wire [$signed(P[1672-:32]) - 1:0] PPN;
			always @(*) begin
				if (_sv2v_0)
					;
				case (WalkerState)
					4'd6, 4'd7: VPN = TranslationVAdr[47:39];
					4'd4, 4'd5: VPN = TranslationVAdr[38:30];
					4'd2, 4'd3: VPN = TranslationVAdr[29:21];
					default: VPN = TranslationVAdr[20:12];
				endcase
			end
			assign PPN = (((WalkerState == 4'd6) | (WalkerState == 4'd7)) | ((SvMode != P[1500-:4]) & ((WalkerState == 4'd4) | (WalkerState == 4'd5))) ? BasePageTablePPN : CurrentPPN);
			assign HPTWReadAdr = {PPN, VPN, 3'b000};
			assign HPTWSize = 3'b011;
		end
		if ($signed(P[4216-:32]) == 32) begin : genblk4
			assign InitialWalkerState = 4'd2;
			assign MegapageMisaligned = |CurrentPPN[9:0];
			assign Misaligned = (WalkerState == 4'd0) & MegapageMisaligned;
		end
		else begin : genblk4
			wire GigapageMisaligned;
			wire TerapageMisaligned;
			assign InitialWalkerState = (SvMode == P[1500-:4] ? 4'd6 : 4'd4);
			assign TerapageMisaligned = |CurrentPPN[26:0];
			assign GigapageMisaligned = |CurrentPPN[17:0];
			assign MegapageMisaligned = |CurrentPPN[8:0];
			assign Misaligned = (((WalkerState == 4'd4) & TerapageMisaligned) | ((WalkerState == 4'd2) & GigapageMisaligned)) | ((WalkerState == 4'd0) & MegapageMisaligned);
		end
	endgenerate
	flopenl_FC78A WalkerStateReg(
		.clk(clk),
		.load(reset | FlushW),
		.en(1'b1),
		.d(NextWalkerState),
		.val(4'd9),
		.q(WalkerState)
	);
	always @(*) begin
		if (_sv2v_0)
			;
		case (WalkerState)
			4'd9:
				if (TLBMissOrUpdateDA)
					NextWalkerState = InitialWalkerState;
				else
					NextWalkerState = 4'd9;
			4'd6: NextWalkerState = 4'd7;
			4'd7:
				if (HPTWFaultM)
					NextWalkerState = 4'd11;
				else if (DCacheBusStallM)
					NextWalkerState = 4'd7;
				else
					NextWalkerState = 4'd4;
			4'd4:
				if (HPTWFaultM)
					NextWalkerState = 4'd11;
				else if ((InitialWalkerState == 4'd4) | ValidNonLeafPTE)
					NextWalkerState = 4'd5;
				else
					NextWalkerState = 4'd8;
			4'd5:
				if (HPTWFaultM)
					NextWalkerState = 4'd11;
				else if (DCacheBusStallM)
					NextWalkerState = 4'd5;
				else
					NextWalkerState = 4'd2;
			4'd2:
				if (HPTWFaultM)
					NextWalkerState = 4'd11;
				else if ((InitialWalkerState == 4'd2) | ValidNonLeafPTE)
					NextWalkerState = 4'd3;
				else
					NextWalkerState = 4'd8;
			4'd3:
				if (HPTWFaultM)
					NextWalkerState = 4'd11;
				else if (DCacheBusStallM)
					NextWalkerState = 4'd3;
				else
					NextWalkerState = 4'd0;
			4'd0:
				if (HPTWFaultM)
					NextWalkerState = 4'd11;
				else if (ValidNonLeafPTE)
					NextWalkerState = 4'd1;
				else
					NextWalkerState = 4'd8;
			4'd1:
				if (HPTWFaultM)
					NextWalkerState = 4'd11;
				else if (DCacheBusStallM)
					NextWalkerState = 4'd1;
				else
					NextWalkerState = 4'd8;
			4'd8:
				if (P[4064] & HPTWUpdateDA)
					NextWalkerState = 4'd10;
				else
					NextWalkerState = 4'd9;
			4'd10:
				if (DCacheBusStallM)
					NextWalkerState = 4'd10;
				else
					NextWalkerState = 4'd8;
			4'd11: NextWalkerState = 4'd9;
			default: NextWalkerState = 4'd9;
		endcase
	end
	assign HPTWFlushW = ((WalkerState == 4'd9) & TLBMissOrUpdateDA) | ((WalkerState != 4'd9) & HPTWFaultM);
	assign SelHPTW = WalkerState != 4'd9;
	assign HPTWStall = ((WalkerState != 4'd9) & (WalkerState != 4'd11)) | ((WalkerState == 4'd9) & TLBMissOrUpdateDA);
	assign SelHPTWAdr = SelHPTW & ~(DTLBWriteM | ITLBWriteF);
	generate
		if ($signed(P[4216-:32]) == 64) begin : genblk5
			assign HPTWAdrExt = {{($signed(P[4216-:32]) + 2) - $signed(P[1640-:32]) {1'b0}}, HPTWAdr};
		end
		else begin : genblk5
			assign HPTWAdrExt = HPTWAdr;
		end
	endgenerate
	mux2 #(.WIDTH(2)) rwmux(
		.d0(MemRWM),
		.d1(HPTWRW),
		.s(SelHPTW),
		.y(PreLSURWM)
	);
	mux2 #(.WIDTH(3)) sizemux(
		.d0(Funct3M),
		.d1(HPTWSize),
		.s(SelHPTW),
		.y(LSUFunct3M)
	);
	mux2 #(.WIDTH(7)) funct7mux(
		.d0(Funct7M),
		.d1(7'b0000000),
		.s(SelHPTW),
		.y(LSUFunct7M)
	);
	mux2 #(.WIDTH(2)) atomicmux(
		.d0(AtomicM),
		.d1(2'b00),
		.s(SelHPTW),
		.y(LSUAtomicM)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]) + 2)) lsupadrmux(
		.d0(IEUAdrExtM),
		.d1(HPTWAdrExt),
		.s(SelHPTWAdr),
		.y(IHAdrM)
	);
	generate
		if (P[4064]) begin : genblk6
			mux2 #(.WIDTH($signed(P[4216-:32]))) lsuwritedatamux(
				.d0(WriteDataM),
				.d1(PTE),
				.s(SelHPTW),
				.y(IHWriteDataM)
			);
		end
		else begin : genblk6
			assign IHWriteDataM = WriteDataM;
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module mmu (
	clk,
	reset,
	SATP_REGW,
	STATUS_MXR,
	STATUS_SUM,
	STATUS_MPRV,
	STATUS_MPP,
	ENVCFG_PBMTE,
	ENVCFG_ADUE,
	PrivilegeModeW,
	DisableTranslation,
	VAdr,
	Size,
	PTE,
	PageTypeWriteVal,
	TLBWrite,
	TLBFlush,
	PhysicalAddress,
	TLBMiss,
	Cacheable,
	Idempotent,
	SelTIM,
	InstrAccessFaultF,
	LoadAccessFaultM,
	StoreAmoAccessFaultM,
	InstrPageFaultF,
	LoadPageFaultM,
	StoreAmoPageFaultM,
	UpdateDA,
	LoadMisalignedFaultM,
	StoreAmoMisalignedFaultM,
	CMOpM,
	AtomicAccessM,
	ExecuteAccessF,
	WriteAccessM,
	ReadAccessM,
	PMPCFG_ARRAY_REGW,
	PMPADDR_ARRAY_REGW
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter TLB_ENTRIES = 8;
	parameter IMMU = 0;
	input wire clk;
	input wire reset;
	input wire [$signed(P[4216-:32]) - 1:0] SATP_REGW;
	input wire STATUS_MXR;
	input wire STATUS_SUM;
	input wire STATUS_MPRV;
	input wire [1:0] STATUS_MPP;
	input wire ENVCFG_PBMTE;
	input wire ENVCFG_ADUE;
	input wire [1:0] PrivilegeModeW;
	input wire DisableTranslation;
	input wire [$signed(P[4216-:32]) + 1:0] VAdr;
	input wire [1:0] Size;
	input wire [$signed(P[4216-:32]) - 1:0] PTE;
	input wire [1:0] PageTypeWriteVal;
	input wire TLBWrite;
	input wire TLBFlush;
	output wire [$signed(P[1640-:32]) - 1:0] PhysicalAddress;
	output wire TLBMiss;
	output wire Cacheable;
	output wire Idempotent;
	output wire SelTIM;
	output wire InstrAccessFaultF;
	output wire LoadAccessFaultM;
	output wire StoreAmoAccessFaultM;
	output wire InstrPageFaultF;
	output wire LoadPageFaultM;
	output wire StoreAmoPageFaultM;
	output wire UpdateDA;
	output wire LoadMisalignedFaultM;
	output wire StoreAmoMisalignedFaultM;
	input wire [3:0] CMOpM;
	input wire AtomicAccessM;
	input wire ExecuteAccessF;
	input wire WriteAccessM;
	input wire ReadAccessM;
	input wire [($signed(P[3728-:32]) * 8) - 1:0] PMPCFG_ARRAY_REGW;
	input wire [(($signed(P[1640-:32]) - 3) >= 0 ? ($signed(P[3728-:32]) * ($signed(P[1640-:32]) - 2)) - 1 : ($signed(P[3728-:32]) * (4 - $signed(P[1640-:32]))) + ($signed(P[1640-:32]) - 4)):(($signed(P[1640-:32]) - 3) >= 0 ? 0 : $signed(P[1640-:32]) - 3)] PMPADDR_ARRAY_REGW;
	wire [$signed(P[1640-:32]) - 1:0] TLBPAdr;
	wire PMAInstrAccessFaultF;
	wire PMPInstrAccessFaultF;
	wire PMALoadAccessFaultM;
	wire PMPLoadAccessFaultM;
	wire PMAStoreAmoAccessFaultM;
	wire PMPStoreAmoAccessFaultM;
	reg DataMisalignedM;
	wire Translate;
	wire TLBPageFault;
	wire ReadNoAmoAccessM;
	wire [1:0] PBMemoryType;
	wire AtomicMisalignedCausesAccessFaultM;
	wire [1:0] EffectivePrivilegeModeW;
	assign EffectivePrivilegeModeW = (IMMU ? PrivilegeModeW : (STATUS_MPRV ? STATUS_MPP : PrivilegeModeW));
	generate
		if (P[4067]) begin : tlb
			wire ReadAccess;
			wire WriteAccess;
			assign ReadAccess = ExecuteAccessF | ReadAccessM;
			assign WriteAccess = WriteAccessM;
			tlb #(
				.P(P),
				.TLB_ENTRIES(TLB_ENTRIES),
				.ITLB(IMMU)
			) tlb(
				.clk(clk),
				.reset(reset),
				.SATP_MODE(SATP_REGW[$signed(P[4216-:32]) - 1:$signed(P[4216-:32]) - $signed(P[1608-:32])]),
				.SATP_ASID(SATP_REGW[($signed(P[1576-:32]) + $signed(P[1544-:32])) - 1:$signed(P[1576-:32])]),
				.VAdr(VAdr[$signed(P[4216-:32]) - 1:0]),
				.STATUS_MXR(STATUS_MXR),
				.STATUS_SUM(STATUS_SUM),
				.STATUS_MPRV(STATUS_MPRV),
				.STATUS_MPP(STATUS_MPP),
				.ENVCFG_PBMTE(ENVCFG_PBMTE),
				.ENVCFG_ADUE(ENVCFG_ADUE),
				.EffectivePrivilegeModeW(EffectivePrivilegeModeW),
				.ReadAccess(ReadAccess),
				.WriteAccess(WriteAccess),
				.CMOpM(CMOpM),
				.DisableTranslation(DisableTranslation),
				.PTE(PTE),
				.PageTypeWriteVal(PageTypeWriteVal),
				.TLBWrite(TLBWrite),
				.TLBFlush(TLBFlush),
				.TLBPAdr(TLBPAdr),
				.TLBMiss(TLBMiss),
				.Translate(Translate),
				.TLBPageFault(TLBPageFault),
				.UpdateDA(UpdateDA),
				.PBMemoryType(PBMemoryType)
			);
		end
		else begin : tlb
			assign Translate = 1'b0;
			assign TLBMiss = 1'b0;
			assign TLBPageFault = 1'b0;
			assign PBMemoryType = 2'b00;
			assign UpdateDA = 1'b0;
			assign TLBPAdr = 1'sb0;
		end
	endgenerate
	mux2 #(.WIDTH($signed(P[1640-:32]) - 12)) addressmux(
		.d0(VAdr[$signed(P[1640-:32]) - 1:12]),
		.d1(TLBPAdr[$signed(P[1640-:32]) - 1:12]),
		.s(Translate),
		.y(PhysicalAddress[$signed(P[1640-:32]) - 1:12])
	);
	assign PhysicalAddress[11:0] = VAdr[11:0];
	pmachecker #(.P(P)) pmachecker(
		.PhysicalAddress(PhysicalAddress),
		.Size(Size),
		.CMOpM(CMOpM),
		.AtomicAccessM(AtomicAccessM),
		.ExecuteAccessF(ExecuteAccessF),
		.WriteAccessM(WriteAccessM),
		.ReadAccessM(ReadAccessM),
		.PBMemoryType(PBMemoryType),
		.Cacheable(Cacheable),
		.Idempotent(Idempotent),
		.SelTIM(SelTIM),
		.PMAInstrAccessFaultF(PMAInstrAccessFaultF),
		.PMALoadAccessFaultM(PMALoadAccessFaultM),
		.PMAStoreAmoAccessFaultM(PMAStoreAmoAccessFaultM)
	);
	generate
		if ($signed(P[3728-:32]) > 0) begin : pmp
			pmpchecker #(.P(P)) pmpchecker(
				.PhysicalAddress(PhysicalAddress),
				.EffectivePrivilegeModeW(EffectivePrivilegeModeW),
				.PMPCFG_ARRAY_REGW(PMPCFG_ARRAY_REGW),
				.PMPADDR_ARRAY_REGW(PMPADDR_ARRAY_REGW),
				.ExecuteAccessF(ExecuteAccessF),
				.WriteAccessM(WriteAccessM),
				.ReadAccessM(ReadAccessM),
				.Size(Size),
				.CMOpM(CMOpM),
				.PMPInstrAccessFaultF(PMPInstrAccessFaultF),
				.PMPLoadAccessFaultM(PMPLoadAccessFaultM),
				.PMPStoreAmoAccessFaultM(PMPStoreAmoAccessFaultM)
			);
		end
		else begin : genblk2
			assign PMPInstrAccessFaultF = 1'b0;
			assign PMPStoreAmoAccessFaultM = 1'b0;
			assign PMPLoadAccessFaultM = 1'b0;
		end
	endgenerate
	assign ReadNoAmoAccessM = ReadAccessM & ~WriteAccessM;
	always @(*) begin
		if (_sv2v_0)
			;
		case (Size)
			2'b00: DataMisalignedM = 1'b0;
			2'b01: DataMisalignedM = VAdr[0];
			2'b10: DataMisalignedM = VAdr[1] | VAdr[0];
			2'b11: DataMisalignedM = |VAdr[2:0];
		endcase
	end
	assign LoadMisalignedFaultM = ((DataMisalignedM & ReadNoAmoAccessM) & ~(P[4059] & Cacheable)) & ~TLBMiss;
	assign StoreAmoMisalignedFaultM = ((DataMisalignedM & WriteAccessM) & ~(P[4059] & Cacheable)) & ~TLBMiss;
	assign AtomicMisalignedCausesAccessFaultM = (DataMisalignedM & AtomicAccessM) & (P[4059] & Cacheable);
	assign InstrAccessFaultF = (PMAInstrAccessFaultF | PMPInstrAccessFaultF) & ~TLBMiss;
	assign LoadAccessFaultM = ((PMALoadAccessFaultM | PMPLoadAccessFaultM) | (AtomicMisalignedCausesAccessFaultM & ReadNoAmoAccessM)) & ~TLBMiss;
	assign StoreAmoAccessFaultM = ((PMAStoreAmoAccessFaultM | PMPStoreAmoAccessFaultM) | (AtomicMisalignedCausesAccessFaultM & WriteAccessM)) & ~TLBMiss;
	assign InstrPageFaultF = TLBPageFault & ExecuteAccessF;
	assign LoadPageFaultM = TLBPageFault & ReadNoAmoAccessM;
	assign StoreAmoPageFaultM = TLBPageFault & (WriteAccessM | (|CMOpM));
	initial _sv2v_0 = 0;
endmodule
module pmachecker (
	PhysicalAddress,
	Size,
	CMOpM,
	AtomicAccessM,
	ExecuteAccessF,
	WriteAccessM,
	ReadAccessM,
	PBMemoryType,
	Cacheable,
	Idempotent,
	SelTIM,
	PMAInstrAccessFaultF,
	PMALoadAccessFaultM,
	PMAStoreAmoAccessFaultM
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[1640-:32]) - 1:0] PhysicalAddress;
	input wire [1:0] Size;
	input wire [3:0] CMOpM;
	input wire AtomicAccessM;
	input wire ExecuteAccessF;
	input wire WriteAccessM;
	input wire ReadAccessM;
	input wire [1:0] PBMemoryType;
	output wire Cacheable;
	output wire Idempotent;
	output wire SelTIM;
	output wire PMAInstrAccessFaultF;
	output wire PMALoadAccessFaultM;
	output wire PMAStoreAmoAccessFaultM;
	wire PMAAccessFault;
	wire AccessRW;
	wire AccessRWXC;
	wire AccessRX;
	wire [11:0] SelRegions;
	wire AtomicAllowed;
	wire CacheableRegion;
	wire IdempotentRegion;
	assign AccessRW = ReadAccessM | WriteAccessM;
	assign AccessRWXC = ((ReadAccessM | WriteAccessM) | ExecuteAccessF) | (|CMOpM);
	assign AccessRX = ReadAccessM | ExecuteAccessF;
	adrdecs #(.P(P)) adrdecs(
		.PhysicalAddress(PhysicalAddress),
		.AccessRW(AccessRW),
		.AccessRX(AccessRX),
		.AccessRWXC(AccessRWXC),
		.Size(Size),
		.SelRegions(SelRegions)
	);
	assign CacheableRegion = (SelRegions[3] | SelRegions[4]) | SelRegions[5];
	assign Cacheable = (PBMemoryType == 2'b00 ? CacheableRegion : 1'b0);
	assign IdempotentRegion = (((SelRegions[1] | SelRegions[2]) | SelRegions[3]) | SelRegions[4]) | SelRegions[5];
	assign Idempotent = (PBMemoryType == 2'b00 ? IdempotentRegion : PBMemoryType == 2'b01);
	assign AtomicAllowed = (SelRegions[1] | SelRegions[3]) | SelRegions[5];
	assign SelTIM = SelRegions[1] | SelRegions[2];
	assign PMAAccessFault = (SelRegions[0] & AccessRWXC) | (AtomicAccessM & ~AtomicAllowed);
	assign PMAInstrAccessFaultF = ExecuteAccessF & PMAAccessFault;
	assign PMALoadAccessFaultM = (ReadAccessM & ~WriteAccessM) & PMAAccessFault;
	assign PMAStoreAmoAccessFaultM = (WriteAccessM | (|CMOpM)) & PMAAccessFault;
endmodule
module pmpadrdec (
	PhysicalAddress,
	Size,
	PMPCfg,
	PMPAdr,
	FirstMatch,
	PAgePMPAdrIn,
	PAgePMPAdrOut,
	Match,
	PMPTop,
	L,
	X,
	W,
	R
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[1640-:32]) - 1:0] PhysicalAddress;
	input wire [1:0] Size;
	input wire [7:0] PMPCfg;
	input wire [$signed(P[1640-:32]) - 3:0] PMPAdr;
	input wire FirstMatch;
	input wire PAgePMPAdrIn;
	output wire PAgePMPAdrOut;
	output wire Match;
	output wire [$signed(P[1640-:32]) - 1:0] PMPTop;
	output wire L;
	output wire X;
	output wire W;
	output wire R;
	localparam TOR = 2'b01;
	localparam NA4 = 2'b10;
	localparam NAPOT = 2'b11;
	wire TORMatch;
	wire NAMatch;
	wire PAltPMPAdr;
	wire [$signed(P[1640-:32]) - 1:0] CurrentAdrFull;
	wire [1:0] AdrMode;
	wire [$signed(P[1640-:32]) - 1:0] PMPTop1;
	wire [$signed(P[1640-:32]) - 1:0] PMPTopTOR;
	wire [$signed(P[1640-:32]) - 1:0] PMPTopNaturallyAligned;
	assign AdrMode = PMPCfg[4:3];
	assign CurrentAdrFull = {PMPAdr, 2'b00};
	assign PAltPMPAdr = {1'b0, PhysicalAddress} < {1'b0, CurrentAdrFull};
	assign PAgePMPAdrOut = ~PAltPMPAdr;
	assign TORMatch = PAgePMPAdrIn & PAltPMPAdr;
	wire [$signed(P[1640-:32]) - 1:0] NAMask;
	wire [$signed(P[1640-:32]) - 1:0] NABase;
	assign NAMask[1:0] = 2'b11;
	assign NAMask[$signed(P[1640-:32]) - 1:2] = (PMPAdr + {{$signed(P[1640-:32]) - 3 {1'b0}}, AdrMode == NAPOT}) ^ PMPAdr;
	assign NABase = {PMPAdr & ~NAMask[$signed(P[1640-:32]) - 1:2], 2'b00};
	assign NAMatch = &((NABase ~^ PhysicalAddress) | NAMask);
	assign Match = (AdrMode == TOR ? TORMatch : ((AdrMode == NA4) | (AdrMode == NAPOT) ? NAMatch : 1'b0));
	assign PMPTopTOR = {PMPAdr - 1, 2'b11};
	assign PMPTopNaturallyAligned = {PMPAdr, 2'b00} | NAMask;
	assign PMPTop1 = (AdrMode == TOR ? PMPTopTOR : PMPTopNaturallyAligned);
	assign PMPTop = (FirstMatch ? PMPTop1 : {$signed(P[1640-:32]) {1'sb0}});
	assign L = PMPCfg[7];
	assign X = PMPCfg[2];
	assign W = PMPCfg[1];
	assign R = PMPCfg[0];
endmodule
module pmpchecker (
	PhysicalAddress,
	EffectivePrivilegeModeW,
	PMPCFG_ARRAY_REGW,
	PMPADDR_ARRAY_REGW,
	ExecuteAccessF,
	WriteAccessM,
	ReadAccessM,
	Size,
	CMOpM,
	PMPInstrAccessFaultF,
	PMPLoadAccessFaultM,
	PMPStoreAmoAccessFaultM
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[1640-:32]) - 1:0] PhysicalAddress;
	input wire [1:0] EffectivePrivilegeModeW;
	input wire [($signed(P[3728-:32]) * 8) - 1:0] PMPCFG_ARRAY_REGW;
	input wire [(($signed(P[1640-:32]) - 3) >= 0 ? ($signed(P[3728-:32]) * ($signed(P[1640-:32]) - 2)) - 1 : ($signed(P[3728-:32]) * (4 - $signed(P[1640-:32]))) + ($signed(P[1640-:32]) - 4)):(($signed(P[1640-:32]) - 3) >= 0 ? 0 : $signed(P[1640-:32]) - 3)] PMPADDR_ARRAY_REGW;
	input wire ExecuteAccessF;
	input wire WriteAccessM;
	input wire ReadAccessM;
	input wire [1:0] Size;
	input wire [3:0] CMOpM;
	output wire PMPInstrAccessFaultF;
	output wire PMPLoadAccessFaultM;
	output wire PMPStoreAmoAccessFaultM;
	wire EnforcePMP;
	wire [$signed(P[3728-:32]) - 1:0] Match;
	wire [$signed(P[3728-:32]) - 1:0] FirstMatch;
	wire [$signed(P[3728-:32]) - 1:0] L;
	wire [$signed(P[3728-:32]) - 1:0] X;
	wire [$signed(P[3728-:32]) - 1:0] W;
	wire [$signed(P[3728-:32]) - 1:0] R;
	wire [$signed(P[3728-:32]) - 1:0] PAgePMPAdr;
	wire [($signed(P[3728-:32]) * $signed(P[1640-:32])) - 1:0] PMPTop;
	wire PMPCMOAccessFault;
	wire PMPCBOMAccessFault;
	wire PMPCBOZAccessFault;
	reg [2:0] SizeBytesMinus1;
	wire MatchingR;
	wire MatchingW;
	wire MatchingX;
	wire MatchingL;
	wire [$signed(P[1640-:32]) - 1:0] MatchingPMPTop;
	wire [$signed(P[1640-:32]) - 1:0] PhysicalAddressTop;
	wire TooBig;
	generate
		if ($signed(P[3728-:32]) > 0) begin : pmp
			pmpadrdec #(.P(P)) pmpadrdecs[$signed(P[3728-:32]) - 1:0](
				.PhysicalAddress(PhysicalAddress),
				.Size(Size),
				.PMPCfg(PMPCFG_ARRAY_REGW),
				.PMPAdr(PMPADDR_ARRAY_REGW),
				.FirstMatch(FirstMatch),
				.PAgePMPAdrIn({PAgePMPAdr[$signed(P[3728-:32]) - 2:0], 1'b1}),
				.PAgePMPAdrOut(PAgePMPAdr),
				.Match(Match),
				.PMPTop(PMPTop),
				.L(L),
				.X(X),
				.W(W),
				.R(R)
			);
		end
	endgenerate
	priorityonehot #(.N($signed(P[3728-:32]))) pmppriority(
		.a(Match),
		.y(FirstMatch)
	);
	assign MatchingR = |(R & FirstMatch) & ~TooBig;
	assign MatchingW = |(W & FirstMatch) & ~TooBig;
	assign MatchingX = |(X & FirstMatch) & ~TooBig;
	assign MatchingL = |(L & FirstMatch);
	or_rows #(
		.ROWS($signed(P[3728-:32])),
		.COLS($signed(P[1640-:32]))
	) PTEOr(
		.a(PMPTop),
		.y(MatchingPMPTop)
	);
	always @(*) begin
		if (_sv2v_0)
			;
		case (Size)
			2'b00: SizeBytesMinus1 = 3'd0;
			2'b01: SizeBytesMinus1 = 3'd1;
			2'b10: SizeBytesMinus1 = 3'd3;
			2'b11: SizeBytesMinus1 = 3'd7;
		endcase
	end
	assign PhysicalAddressTop = PhysicalAddress + {{$signed(P[1640-:32]) - 3 {1'b0}}, SizeBytesMinus1};
	assign TooBig = PhysicalAddressTop > MatchingPMPTop;
	assign EnforcePMP = (EffectivePrivilegeModeW != P[1742-:2]) | MatchingL;
	assign PMPCBOMAccessFault = (EnforcePMP & |CMOpM[2:0]) & ~MatchingR;
	assign PMPCBOZAccessFault = (EnforcePMP & CMOpM[3]) & ~MatchingW;
	assign PMPCMOAccessFault = PMPCBOZAccessFault | PMPCBOMAccessFault;
	assign PMPInstrAccessFaultF = (EnforcePMP & ExecuteAccessF) & ~MatchingX;
	assign PMPStoreAmoAccessFaultM = ((EnforcePMP & WriteAccessM) & ~MatchingW) | PMPCMOAccessFault;
	assign PMPLoadAccessFaultM = ((EnforcePMP & ReadAccessM) & ~WriteAccessM) & ~MatchingR;
	initial _sv2v_0 = 0;
endmodule
module csr (
	clk,
	reset,
	FlushM,
	FlushW,
	StallE,
	StallM,
	StallW,
	InstrM,
	InstrOrigM,
	PCM,
	SrcAM,
	IEUAdrxTvalM,
	CSRReadM,
	CSRWriteM,
	TrapM,
	mretM,
	sretM,
	InterruptM,
	ExceptionM,
	MTimerInt,
	MExtInt,
	SExtInt,
	MSwInt,
	MTIME_CLINT,
	InstrValidM,
	FRegWriteM,
	SetFflagsM,
	NextPrivilegeModeM,
	PrivilegeModeW,
	CauseM,
	SelHPTW,
	LoadStallD,
	StoreStallD,
	ICacheStallF,
	DCacheStallM,
	BPDirWrongM,
	BTAWrongM,
	RASPredPCWrongM,
	IClassWrongM,
	BPWrongM,
	IClassM,
	DCacheMiss,
	DCacheAccess,
	ICacheMiss,
	ICacheAccess,
	sfencevmaM,
	InvalidateICacheM,
	DivBusyE,
	FDivBusyE,
	STATUS_MPP,
	STATUS_SPP,
	STATUS_TSR,
	STATUS_TVM,
	MEDELEG_REGW,
	SATP_REGW,
	MIP_REGW,
	MIE_REGW,
	MIDELEG_REGW,
	STATUS_MIE,
	STATUS_SIE,
	STATUS_MXR,
	STATUS_SUM,
	STATUS_MPRV,
	STATUS_TW,
	STATUS_FS,
	PMPCFG_ARRAY_REGW,
	PMPADDR_ARRAY_REGW,
	FRM_REGW,
	ENVCFG_CBE,
	ENVCFG_PBMTE,
	ENVCFG_ADUE,
	EPCM,
	TrapVectorM,
	CSRReadValW,
	IllegalCSRAccessM,
	BigEndianM
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire FlushM;
	input wire FlushW;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire [31:0] InstrM;
	input wire [31:0] InstrOrigM;
	input wire [$signed(P[4216-:32]) - 1:0] PCM;
	input wire [$signed(P[4216-:32]) - 1:0] SrcAM;
	input wire [$signed(P[4216-:32]) - 1:0] IEUAdrxTvalM;
	input wire CSRReadM;
	input wire CSRWriteM;
	input wire TrapM;
	input wire mretM;
	input wire sretM;
	input wire InterruptM;
	input wire ExceptionM;
	input wire MTimerInt;
	input wire MExtInt;
	input wire SExtInt;
	input wire MSwInt;
	input wire [63:0] MTIME_CLINT;
	input wire InstrValidM;
	input wire FRegWriteM;
	input wire [4:0] SetFflagsM;
	input wire [1:0] NextPrivilegeModeM;
	input wire [1:0] PrivilegeModeW;
	input wire [3:0] CauseM;
	input wire SelHPTW;
	input wire LoadStallD;
	input wire StoreStallD;
	input wire ICacheStallF;
	input wire DCacheStallM;
	input wire BPDirWrongM;
	input wire BTAWrongM;
	input wire RASPredPCWrongM;
	input wire IClassWrongM;
	input wire BPWrongM;
	input wire [3:0] IClassM;
	input wire DCacheMiss;
	input wire DCacheAccess;
	input wire ICacheMiss;
	input wire ICacheAccess;
	input wire sfencevmaM;
	input wire InvalidateICacheM;
	input wire DivBusyE;
	input wire FDivBusyE;
	output wire [1:0] STATUS_MPP;
	output wire STATUS_SPP;
	output wire STATUS_TSR;
	output wire STATUS_TVM;
	output wire [15:0] MEDELEG_REGW;
	output wire [$signed(P[4216-:32]) - 1:0] SATP_REGW;
	output wire [11:0] MIP_REGW;
	output wire [11:0] MIE_REGW;
	output wire [11:0] MIDELEG_REGW;
	output wire STATUS_MIE;
	output wire STATUS_SIE;
	output wire STATUS_MXR;
	output wire STATUS_SUM;
	output wire STATUS_MPRV;
	output wire STATUS_TW;
	output wire [1:0] STATUS_FS;
	output wire [($signed(P[3728-:32]) * 8) - 1:0] PMPCFG_ARRAY_REGW;
	output wire [(($signed(P[1640-:32]) - 3) >= 0 ? ($signed(P[3728-:32]) * ($signed(P[1640-:32]) - 2)) - 1 : ($signed(P[3728-:32]) * (4 - $signed(P[1640-:32]))) + ($signed(P[1640-:32]) - 4)):(($signed(P[1640-:32]) - 3) >= 0 ? 0 : $signed(P[1640-:32]) - 3)] PMPADDR_ARRAY_REGW;
	output wire [2:0] FRM_REGW;
	output wire [3:0] ENVCFG_CBE;
	output wire ENVCFG_PBMTE;
	output wire ENVCFG_ADUE;
	output wire [$signed(P[4216-:32]) - 1:0] EPCM;
	output wire [$signed(P[4216-:32]) - 1:0] TrapVectorM;
	output wire [$signed(P[4216-:32]) - 1:0] CSRReadValW;
	output wire IllegalCSRAccessM;
	output wire BigEndianM;
	localparam MIP = 12'h344;
	localparam SIP = 12'h144;
	wire [$signed(P[4216-:32]) - 1:0] CSRMReadValM;
	wire [$signed(P[4216-:32]) - 1:0] CSRSReadValM;
	wire [$signed(P[4216-:32]) - 1:0] CSRUReadValM;
	wire [$signed(P[4216-:32]) - 1:0] CSRCReadValM;
	wire [$signed(P[4216-:32]) - 1:0] CSRReadValM;
	reg [$signed(P[4216-:32]) - 1:0] CSRSrcM;
	reg [$signed(P[4216-:32]) - 1:0] CSRRWM;
	reg [$signed(P[4216-:32]) - 1:0] CSRRSM;
	reg [$signed(P[4216-:32]) - 1:0] CSRRCM;
	reg [$signed(P[4216-:32]) - 1:0] CSRWriteValM;
	wire [$signed(P[4216-:32]) - 1:0] MSTATUS_REGW;
	wire [$signed(P[4216-:32]) - 1:0] SSTATUS_REGW;
	wire [$signed(P[4216-:32]) - 1:0] MSTATUSH_REGW;
	wire [$signed(P[4216-:32]) - 1:0] STVEC_REGW;
	wire [$signed(P[4216-:32]) - 1:0] MTVEC_REGW;
	wire [$signed(P[4216-:32]) - 1:0] MEPC_REGW;
	wire [$signed(P[4216-:32]) - 1:0] SEPC_REGW;
	wire [31:0] MCOUNTINHIBIT_REGW;
	wire [31:0] MCOUNTEREN_REGW;
	wire [31:0] SCOUNTEREN_REGW;
	wire WriteMSTATUSM;
	wire WriteMSTATUSHM;
	wire WriteSSTATUSM;
	wire CSRMWriteM;
	wire CSRSWriteM;
	wire CSRUWriteM;
	wire UngatedCSRMWriteM;
	wire WriteFRMM;
	wire SetOrWriteFFLAGSM;
	wire [$signed(P[4216-:32]) - 1:0] UnalignedNextEPCM;
	wire [$signed(P[4216-:32]) - 1:0] NextEPCM;
	wire [$signed(P[4216-:32]) - 1:0] NextMtvalM;
	wire [4:0] NextCauseM;
	wire [11:0] CSRAdrM;
	wire IllegalCSRCAccessM;
	wire IllegalCSRMAccessM;
	wire IllegalCSRSAccessM;
	wire IllegalCSRUAccessM;
	wire InsufficientCSRPrivilegeM;
	wire IllegalCSRMWriteReadonlyM;
	reg [$signed(P[4216-:32]) - 1:0] CSRReadVal2M;
	wire [11:0] MIP_REGW_writeable;
	wire [$signed(P[4216-:32]) - 1:0] TVecM;
	reg [$signed(P[4216-:32]) - 1:0] NextFaultMtvalM;
	wire MTrapM;
	wire STrapM;
	wire SelMtvecM;
	wire [$signed(P[4216-:32]) - 1:0] TVecAlignedM;
	wire InstrValidNotFlushedM;
	wire STimerInt;
	wire [63:0] MENVCFG_REGW;
	wire [$signed(P[4216-:32]) - 1:0] SENVCFG_REGW;
	wire ENVCFG_STCE;
	wire ENVCFG_FIOM;
	assign InstrValidNotFlushedM = (InstrValidM & ~StallW) & ~FlushW;
	always @(*) begin
		if (_sv2v_0)
			;
		if (InterruptM)
			NextFaultMtvalM = 1'sb0;
		else
			case (CauseM)
				12, 1, 3: NextFaultMtvalM = PCM;
				2: NextFaultMtvalM = {{$signed(P[4216-:32]) - 32 {1'b0}}, InstrOrigM};
				0, 4, 6, 13, 15, 5, 7: NextFaultMtvalM = IEUAdrxTvalM;
				default: NextFaultMtvalM = 1'sb0;
			endcase
	end
	assign SelMtvecM = NextPrivilegeModeM == P[1742-:2];
	mux2 #(.WIDTH($signed(P[4216-:32]))) tvecmux(
		.d0(STVEC_REGW),
		.d1(MTVEC_REGW),
		.s(SelMtvecM),
		.y(TVecM)
	);
	assign TVecAlignedM = {TVecM[$signed(P[4216-:32]) - 1:2], 2'b00};
	generate
		if (P[4066]) begin : vec
			wire VectoredM;
			wire [$signed(P[4216-:32]) - 1:0] TVecPlusCauseM;
			assign VectoredM = InterruptM & (TVecM[1:0] == 2'b01);
			assign TVecPlusCauseM = {TVecAlignedM[$signed(P[4216-:32]) - 1:6], CauseM, 2'b00};
			mux2 #(.WIDTH($signed(P[4216-:32]))) trapvecmux(
				.d0(TVecAlignedM),
				.d1(TVecPlusCauseM),
				.s(VectoredM),
				.y(TrapVectorM)
			);
		end
		else begin : genblk1
			assign TrapVectorM = TVecAlignedM;
		end
	endgenerate
	mux2 #(.WIDTH($signed(P[4216-:32]))) epcmux(
		.d0(SEPC_REGW),
		.d1(MEPC_REGW),
		.s(mretM),
		.y(EPCM)
	);
	always @(*) begin
		if (_sv2v_0)
			;
		CSRSrcM = (InstrM[14] ? {{$signed(P[4216-:32]) - 5 {1'b0}}, InstrM[19:15]} : SrcAM);
		if ((CSRAdrM == MIP) | (CSRAdrM == SIP))
			CSRReadVal2M = {{$signed(P[4216-:32]) - 12 {1'b0}}, MIP_REGW_writeable};
		else
			CSRReadVal2M = CSRReadValM;
		CSRRWM = CSRSrcM;
		CSRRSM = CSRReadVal2M | CSRSrcM;
		CSRRCM = CSRReadVal2M & ~CSRSrcM;
		case (InstrM[13:12])
			2'b01: CSRWriteValM = CSRRWM;
			2'b10: CSRWriteValM = CSRRSM;
			2'b11: CSRWriteValM = CSRRCM;
			default: CSRWriteValM = CSRReadValM;
		endcase
	end
	assign CSRAdrM = InstrM[31:20];
	assign UnalignedNextEPCM = (TrapM ? PCM : CSRWriteValM);
	assign NextEPCM = (P[1754] ? {UnalignedNextEPCM[$signed(P[4216-:32]) - 1:1], 1'b0} : {UnalignedNextEPCM[$signed(P[4216-:32]) - 1:2], 2'b00});
	assign NextCauseM = (TrapM ? {InterruptM, CauseM} : {CSRWriteValM[$signed(P[4216-:32]) - 1], CSRWriteValM[3:0]});
	assign NextMtvalM = (TrapM ? NextFaultMtvalM : CSRWriteValM);
	assign UngatedCSRMWriteM = CSRWriteM & (PrivilegeModeW == P[1742-:2]);
	assign CSRMWriteM = UngatedCSRMWriteM & InstrValidNotFlushedM;
	assign CSRSWriteM = (CSRWriteM & |PrivilegeModeW) & InstrValidNotFlushedM;
	assign CSRUWriteM = CSRWriteM & InstrValidNotFlushedM;
	assign MTrapM = TrapM & (NextPrivilegeModeM == P[1742-:2]);
	assign STrapM = (TrapM & (NextPrivilegeModeM == P[1740-:2])) & P[1487];
	csri #(.P(P)) csri(
		.clk(clk),
		.reset(reset),
		.CSRMWriteM(CSRMWriteM),
		.CSRSWriteM(CSRSWriteM),
		.CSRWriteValM(CSRWriteValM),
		.CSRAdrM(CSRAdrM),
		.MExtInt(MExtInt),
		.SExtInt(SExtInt),
		.MTimerInt(MTimerInt),
		.STimerInt(STimerInt),
		.MSwInt(MSwInt),
		.MIDELEG_REGW(MIDELEG_REGW),
		.ENVCFG_STCE(ENVCFG_STCE),
		.MIP_REGW(MIP_REGW),
		.MIE_REGW(MIE_REGW),
		.MIP_REGW_writeable(MIP_REGW_writeable)
	);
	csrsr #(.P(P)) csrsr(
		.clk(clk),
		.reset(reset),
		.StallW(StallW),
		.WriteMSTATUSM(WriteMSTATUSM),
		.WriteMSTATUSHM(WriteMSTATUSHM),
		.WriteSSTATUSM(WriteSSTATUSM),
		.TrapM(TrapM),
		.FRegWriteM(FRegWriteM),
		.NextPrivilegeModeM(NextPrivilegeModeM),
		.PrivilegeModeW(PrivilegeModeW),
		.mretM(mretM),
		.sretM(sretM),
		.WriteFRMM(WriteFRMM),
		.SetOrWriteFFLAGSM(SetOrWriteFFLAGSM),
		.CSRWriteValM(CSRWriteValM),
		.SelHPTW(SelHPTW),
		.MSTATUS_REGW(MSTATUS_REGW),
		.SSTATUS_REGW(SSTATUS_REGW),
		.MSTATUSH_REGW(MSTATUSH_REGW),
		.STATUS_MPP(STATUS_MPP),
		.STATUS_SPP(STATUS_SPP),
		.STATUS_TSR(STATUS_TSR),
		.STATUS_TW(STATUS_TW),
		.STATUS_MIE(STATUS_MIE),
		.STATUS_SIE(STATUS_SIE),
		.STATUS_MXR(STATUS_MXR),
		.STATUS_SUM(STATUS_SUM),
		.STATUS_MPRV(STATUS_MPRV),
		.STATUS_TVM(STATUS_TVM),
		.STATUS_FS(STATUS_FS),
		.BigEndianM(BigEndianM)
	);
	csrm #(.P(P)) csrm(
		.clk(clk),
		.reset(reset),
		.UngatedCSRMWriteM(UngatedCSRMWriteM),
		.CSRMWriteM(CSRMWriteM),
		.MTrapM(MTrapM),
		.CSRAdrM(CSRAdrM),
		.NextEPCM(NextEPCM),
		.NextCauseM(NextCauseM),
		.NextMtvalM(NextMtvalM),
		.MSTATUS_REGW(MSTATUS_REGW),
		.MSTATUSH_REGW(MSTATUSH_REGW),
		.CSRWriteValM(CSRWriteValM),
		.CSRMReadValM(CSRMReadValM),
		.MTVEC_REGW(MTVEC_REGW),
		.MEPC_REGW(MEPC_REGW),
		.MCOUNTEREN_REGW(MCOUNTEREN_REGW),
		.MCOUNTINHIBIT_REGW(MCOUNTINHIBIT_REGW),
		.MEDELEG_REGW(MEDELEG_REGW),
		.MIDELEG_REGW(MIDELEG_REGW),
		.PMPCFG_ARRAY_REGW(PMPCFG_ARRAY_REGW),
		.PMPADDR_ARRAY_REGW(PMPADDR_ARRAY_REGW),
		.MIP_REGW(MIP_REGW),
		.MIE_REGW(MIE_REGW),
		.WriteMSTATUSM(WriteMSTATUSM),
		.WriteMSTATUSHM(WriteMSTATUSHM),
		.IllegalCSRMAccessM(IllegalCSRMAccessM),
		.IllegalCSRMWriteReadonlyM(IllegalCSRMWriteReadonlyM),
		.MENVCFG_REGW(MENVCFG_REGW)
	);
	generate
		if (P[1487]) begin : csrs
			wire STCE;
			assign STCE = P[4068] & ((PrivilegeModeW == P[1742-:2]) | (MCOUNTEREN_REGW[1] & ENVCFG_STCE));
			csrs #(.P(P)) csrs(
				.clk(clk),
				.reset(reset),
				.CSRSWriteM(CSRSWriteM),
				.STrapM(STrapM),
				.CSRAdrM(CSRAdrM),
				.NextEPCM(NextEPCM),
				.NextCauseM(NextCauseM),
				.NextMtvalM(NextMtvalM),
				.SSTATUS_REGW(SSTATUS_REGW),
				.STATUS_TVM(STATUS_TVM),
				.CSRWriteValM(CSRWriteValM),
				.PrivilegeModeW(PrivilegeModeW),
				.CSRSReadValM(CSRSReadValM),
				.STVEC_REGW(STVEC_REGW),
				.SEPC_REGW(SEPC_REGW),
				.SCOUNTEREN_REGW(SCOUNTEREN_REGW),
				.SATP_REGW(SATP_REGW),
				.MIP_REGW(MIP_REGW),
				.MIE_REGW(MIE_REGW),
				.MIDELEG_REGW(MIDELEG_REGW),
				.MTIME_CLINT(MTIME_CLINT),
				.STCE(STCE),
				.WriteSSTATUSM(WriteSSTATUSM),
				.IllegalCSRSAccessM(IllegalCSRSAccessM),
				.STimerInt(STimerInt),
				.SENVCFG_REGW(SENVCFG_REGW)
			);
		end
		else begin : genblk2
			assign WriteSSTATUSM = 1'b0;
			assign CSRSReadValM = 1'sb0;
			assign SEPC_REGW = 1'sb0;
			assign STVEC_REGW = 1'sb0;
			assign SCOUNTEREN_REGW = 1'sb0;
			assign SATP_REGW = 1'sb0;
			assign IllegalCSRSAccessM = 1'b1;
			assign STimerInt = 1'sb0;
			assign SENVCFG_REGW = 1'sb0;
		end
		if (P[1491]) begin : csru
			csru #(.P(P)) csru(
				.clk(clk),
				.reset(reset),
				.InstrValidNotFlushedM(InstrValidNotFlushedM),
				.CSRUWriteM(CSRUWriteM),
				.CSRAdrM(CSRAdrM),
				.CSRWriteValM(CSRWriteValM),
				.STATUS_FS(STATUS_FS),
				.CSRUReadValM(CSRUReadValM),
				.SetFflagsM(SetFflagsM),
				.FRM_REGW(FRM_REGW),
				.WriteFRMM(WriteFRMM),
				.SetOrWriteFFLAGSM(SetOrWriteFFLAGSM),
				.IllegalCSRUAccessM(IllegalCSRUAccessM)
			);
		end
		else begin : genblk3
			assign FRM_REGW = 1'sb0;
			assign CSRUReadValM = 1'sb0;
			assign IllegalCSRUAccessM = 1'b1;
			assign WriteFRMM = 1'b0;
			assign SetOrWriteFFLAGSM = 1'b0;
		end
		if (P[4072]) begin : counters
			csrc #(.P(P)) counters(
				.clk(clk),
				.reset(reset),
				.StallE(StallE),
				.StallM(StallM),
				.FlushM(FlushM),
				.InstrValidNotFlushedM(InstrValidNotFlushedM),
				.LoadStallD(LoadStallD),
				.StoreStallD(StoreStallD),
				.CSRWriteM(CSRWriteM),
				.CSRMWriteM(CSRMWriteM),
				.BPDirWrongM(BPDirWrongM),
				.BTAWrongM(BTAWrongM),
				.RASPredPCWrongM(RASPredPCWrongM),
				.IClassWrongM(IClassWrongM),
				.BPWrongM(BPWrongM),
				.IClassM(IClassM),
				.DCacheMiss(DCacheMiss),
				.DCacheAccess(DCacheAccess),
				.ICacheMiss(ICacheMiss),
				.ICacheAccess(ICacheAccess),
				.sfencevmaM(sfencevmaM),
				.InterruptM(InterruptM),
				.ExceptionM(ExceptionM),
				.InvalidateICacheM(InvalidateICacheM),
				.ICacheStallF(ICacheStallF),
				.DCacheStallM(DCacheStallM),
				.DivBusyE(DivBusyE),
				.FDivBusyE(FDivBusyE),
				.CSRAdrM(CSRAdrM),
				.PrivilegeModeW(PrivilegeModeW),
				.CSRWriteValM(CSRWriteValM),
				.MCOUNTINHIBIT_REGW(MCOUNTINHIBIT_REGW),
				.MCOUNTEREN_REGW(MCOUNTEREN_REGW),
				.SCOUNTEREN_REGW(SCOUNTEREN_REGW),
				.MTIME_CLINT(MTIME_CLINT),
				.CSRCReadValM(CSRCReadValM),
				.IllegalCSRCAccessM(IllegalCSRCAccessM)
			);
		end
		else begin : genblk4
			assign CSRCReadValM = 1'sb0;
			assign IllegalCSRCAccessM = 1'b1;
		end
	endgenerate
	assign ENVCFG_STCE = MENVCFG_REGW[63];
	assign ENVCFG_PBMTE = MENVCFG_REGW[62];
	assign ENVCFG_ADUE = MENVCFG_REGW[61];
	assign ENVCFG_CBE = (PrivilegeModeW == P[1742-:2] ? 4'b1111 : ((PrivilegeModeW == P[1740-:2]) | !P[1487] ? MENVCFG_REGW[7:4] : MENVCFG_REGW[7:4] & SENVCFG_REGW[7:4]));
	assign ENVCFG_FIOM = (PrivilegeModeW == P[1742-:2] ? 1'b1 : ((PrivilegeModeW == P[1740-:2]) | !P[1487] ? MENVCFG_REGW[0] : MENVCFG_REGW[0] & SENVCFG_REGW[0]));
	assign CSRReadValM = ((CSRUReadValM | CSRSReadValM) | CSRMReadValM) | CSRCReadValM;
	flopenrc #(.WIDTH($signed(P[4216-:32]))) CSRValWReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(CSRReadValM),
		.q(CSRReadValW)
	);
	assign InsufficientCSRPrivilegeM = ((CSRAdrM[9:8] == 2'b11) & (PrivilegeModeW != P[1742-:2])) | ((CSRAdrM[9:8] == 2'b01) & (PrivilegeModeW == P[1738-:2]));
	assign IllegalCSRAccessM = (((((IllegalCSRCAccessM & IllegalCSRMAccessM) & IllegalCSRSAccessM) & IllegalCSRUAccessM) | InsufficientCSRPrivilegeM) & CSRReadM) | IllegalCSRMWriteReadonlyM;
	initial _sv2v_0 = 0;
endmodule
module csrc (
	clk,
	reset,
	StallE,
	StallM,
	FlushM,
	InstrValidNotFlushedM,
	LoadStallD,
	StoreStallD,
	CSRMWriteM,
	CSRWriteM,
	BPDirWrongM,
	BTAWrongM,
	RASPredPCWrongM,
	IClassWrongM,
	BPWrongM,
	IClassM,
	DCacheMiss,
	DCacheAccess,
	ICacheMiss,
	ICacheAccess,
	ICacheStallF,
	DCacheStallM,
	sfencevmaM,
	InterruptM,
	ExceptionM,
	InvalidateICacheM,
	DivBusyE,
	FDivBusyE,
	CSRAdrM,
	PrivilegeModeW,
	CSRWriteValM,
	MCOUNTINHIBIT_REGW,
	MCOUNTEREN_REGW,
	SCOUNTEREN_REGW,
	MTIME_CLINT,
	CSRCReadValM,
	IllegalCSRCAccessM
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallE;
	input wire StallM;
	input wire FlushM;
	input wire InstrValidNotFlushedM;
	input wire LoadStallD;
	input wire StoreStallD;
	input wire CSRMWriteM;
	input wire CSRWriteM;
	input wire BPDirWrongM;
	input wire BTAWrongM;
	input wire RASPredPCWrongM;
	input wire IClassWrongM;
	input wire BPWrongM;
	input wire [3:0] IClassM;
	input wire DCacheMiss;
	input wire DCacheAccess;
	input wire ICacheMiss;
	input wire ICacheAccess;
	input wire ICacheStallF;
	input wire DCacheStallM;
	input wire sfencevmaM;
	input wire InterruptM;
	input wire ExceptionM;
	input wire InvalidateICacheM;
	input wire DivBusyE;
	input wire FDivBusyE;
	input wire [11:0] CSRAdrM;
	input wire [1:0] PrivilegeModeW;
	input wire [$signed(P[4216-:32]) - 1:0] CSRWriteValM;
	input wire [31:0] MCOUNTINHIBIT_REGW;
	input wire [31:0] MCOUNTEREN_REGW;
	input wire [31:0] SCOUNTEREN_REGW;
	input wire [63:0] MTIME_CLINT;
	output reg [$signed(P[4216-:32]) - 1:0] CSRCReadValM;
	output reg IllegalCSRCAccessM;
	localparam MHPMCOUNTERBASE = 12'hb00;
	localparam MTIME = 12'hb01;
	localparam MHPMCOUNTERHBASE = 12'hb80;
	localparam MTIMEH = 12'hb81;
	localparam MHPMEVENTBASE = 12'h323;
	localparam MHPMEVENTLAST = 12'h33f;
	localparam HPMCOUNTERBASE = 12'hc00;
	localparam HPMCOUNTERHBASE = 12'hc80;
	localparam TIME = 12'hc01;
	localparam TIMEH = 12'hc81;
	wire [4:0] CounterNumM;
	reg [$signed(P[4216-:32]) - 1:0] HPMCOUNTER_REGW [P[4084-:12] - 1:0];
	reg [$signed(P[4216-:32]) - 1:0] HPMCOUNTERH_REGW [P[4084-:12] - 1:0];
	wire LoadStallE;
	wire LoadStallM;
	wire StoreStallE;
	wire StoreStallM;
	wire [P[4084-:12] - 1:0] WriteHPMCOUNTERM;
	wire [P[4084-:12] - 1:0] CounterEvent;
	wire [63:0] HPMCOUNTERPlusM [P[4084-:12] - 1:0];
	wire [$signed(P[4216-:32]) - 1:0] NextHPMCOUNTERM [P[4084-:12] - 1:0];
	genvar _gv_i_4;
	flopenrc #(.WIDTH(1)) LoadStallEReg(
		.clk(clk),
		.reset(reset),
		.clear(1'b0),
		.en(~StallE),
		.d(LoadStallD),
		.q(LoadStallE)
	);
	flopenrc #(.WIDTH(1)) LoadStallMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(LoadStallE),
		.q(LoadStallM)
	);
	flopenrc #(.WIDTH(1)) StoreStallEReg(
		.clk(clk),
		.reset(reset),
		.clear(1'b0),
		.en(~StallE),
		.d(StoreStallD),
		.q(StoreStallE)
	);
	flopenrc #(.WIDTH(1)) StoreStallMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(StoreStallE),
		.q(StoreStallM)
	);
	assign CounterEvent[0] = 1'b1;
	assign CounterEvent[1] = 1'b0;
	assign CounterEvent[2] = InstrValidNotFlushedM;
	generate
		if (P[4071]) begin : cevent
			assign CounterEvent[3] = IClassM[0] & InstrValidNotFlushedM;
			assign CounterEvent[4] = (IClassM[1] & ~IClassM[2]) & InstrValidNotFlushedM;
			assign CounterEvent[5] = IClassM[2] & InstrValidNotFlushedM;
			assign CounterEvent[6] = BPWrongM & InstrValidNotFlushedM;
			assign CounterEvent[7] = BPDirWrongM & InstrValidNotFlushedM;
			assign CounterEvent[8] = BTAWrongM & InstrValidNotFlushedM;
			assign CounterEvent[9] = RASPredPCWrongM & InstrValidNotFlushedM;
			assign CounterEvent[10] = IClassWrongM & InstrValidNotFlushedM;
			assign CounterEvent[11] = LoadStallM;
			assign CounterEvent[12] = StoreStallM;
			assign CounterEvent[13] = DCacheAccess;
			assign CounterEvent[14] = DCacheMiss;
			assign CounterEvent[15] = DCacheStallM;
			assign CounterEvent[16] = ICacheAccess;
			assign CounterEvent[17] = ICacheMiss;
			assign CounterEvent[18] = ICacheStallF;
			assign CounterEvent[19] = CSRWriteM & InstrValidNotFlushedM;
			assign CounterEvent[20] = InvalidateICacheM & InstrValidNotFlushedM;
			assign CounterEvent[21] = sfencevmaM & InstrValidNotFlushedM;
			assign CounterEvent[22] = InterruptM;
			assign CounterEvent[23] = ExceptionM;
			assign CounterEvent[24] = DivBusyE | FDivBusyE;
			assign CounterEvent[P[4084-:12] - 1:25] = 1'sb0;
		end
		else begin : cevent
			assign CounterEvent[P[4084-:12] - 1:3] = 1'sb0;
		end
		for (_gv_i_4 = 0; $unsigned(_gv_i_4) < P[4084-:12]; _gv_i_4 = _gv_i_4 + 1) begin : cntr
			localparam i = _gv_i_4;
			assign WriteHPMCOUNTERM[i] = CSRMWriteM & (CSRAdrM == (MHPMCOUNTERBASE + i));
			assign NextHPMCOUNTERM[i][$signed(P[4216-:32]) - 1:0] = (WriteHPMCOUNTERM[i] ? CSRWriteValM : HPMCOUNTERPlusM[i][$signed(P[4216-:32]) - 1:0]);
			always @(posedge clk)
				if (reset)
					HPMCOUNTER_REGW[i][$signed(P[4216-:32]) - 1:0] <= 1'sb0;
				else
					HPMCOUNTER_REGW[i][$signed(P[4216-:32]) - 1:0] <= NextHPMCOUNTERM[i];
			if ($signed(P[4216-:32]) == 32) begin : genblk1
				wire [P[4084-:12] - 1:0] WriteHPMCOUNTERHM;
				wire [$signed(P[4216-:32]) - 1:0] NextHPMCOUNTERHM [P[4084-:12] - 1:0];
				assign HPMCOUNTERPlusM[i] = {HPMCOUNTERH_REGW[i], HPMCOUNTER_REGW[i]} + {63'b000000000000000000000000000000000000000000000000000000000000000, CounterEvent[i] & ~MCOUNTINHIBIT_REGW[i]};
				assign WriteHPMCOUNTERHM[i] = CSRMWriteM & (CSRAdrM == (MHPMCOUNTERHBASE + i));
				assign NextHPMCOUNTERHM[i] = (WriteHPMCOUNTERHM[i] ? CSRWriteValM : HPMCOUNTERPlusM[i][63:32]);
				always @(posedge clk)
					if (reset)
						HPMCOUNTERH_REGW[i][$signed(P[4216-:32]) - 1:0] <= 1'sb0;
					else
						HPMCOUNTERH_REGW[i][$signed(P[4216-:32]) - 1:0] <= NextHPMCOUNTERHM[i];
			end
			else begin : genblk1
				assign HPMCOUNTERPlusM[i] = HPMCOUNTER_REGW[i] + {63'b000000000000000000000000000000000000000000000000000000000000000, CounterEvent[i] & ~MCOUNTINHIBIT_REGW[i]};
				wire [$signed(P[4216-:32]):1] sv2v_tmp_20CDA;
				assign sv2v_tmp_20CDA = 1'sb0;
				always @(*) HPMCOUNTERH_REGW[i] = sv2v_tmp_20CDA;
			end
		end
	endgenerate
	assign CounterNumM = CSRAdrM[4:0];
	always @(*) begin
		if (_sv2v_0)
			;
		if ((PrivilegeModeW == P[1742-:2]) | (MCOUNTEREN_REGW[CounterNumM] & ((!P[1487] | (PrivilegeModeW == P[1740-:2])) | SCOUNTEREN_REGW[CounterNumM]))) begin
			IllegalCSRCAccessM = 1'b0;
			if ((CSRAdrM >= MHPMEVENTBASE) & (CSRAdrM <= MHPMEVENTLAST))
				CSRCReadValM = 1'sb0;
			else if ($signed(P[4216-:32]) == 64) begin
				if ((CSRAdrM == TIME) & ~CSRWriteM)
					CSRCReadValM = MTIME_CLINT;
				else if (((CSRAdrM >= MHPMCOUNTERBASE) & (CSRAdrM < (MHPMCOUNTERBASE + P[4084-:12]))) & (CSRAdrM != MTIME))
					CSRCReadValM = HPMCOUNTER_REGW[CounterNumM];
				else if (((CSRAdrM >= HPMCOUNTERBASE) & (CSRAdrM < (HPMCOUNTERBASE + P[4084-:12]))) & ~CSRWriteM)
					CSRCReadValM = HPMCOUNTER_REGW[CounterNumM];
				else begin
					CSRCReadValM = 1'sb0;
					IllegalCSRCAccessM = 1'b1;
				end
			end
			else if ((CSRAdrM == TIME) & ~CSRWriteM)
				CSRCReadValM = MTIME_CLINT[31:0];
			else if ((CSRAdrM == TIMEH) & ~CSRWriteM)
				CSRCReadValM = MTIME_CLINT[63:32];
			else if (((CSRAdrM >= MHPMCOUNTERBASE) & (CSRAdrM < (MHPMCOUNTERBASE + P[4084-:12]))) & (CSRAdrM != MTIME))
				CSRCReadValM = HPMCOUNTER_REGW[CounterNumM];
			else if (((CSRAdrM >= HPMCOUNTERBASE) & (CSRAdrM < (HPMCOUNTERBASE + P[4084-:12]))) & ~CSRWriteM)
				CSRCReadValM = HPMCOUNTER_REGW[CounterNumM];
			else if (((CSRAdrM >= MHPMCOUNTERHBASE) & (CSRAdrM < (MHPMCOUNTERHBASE + P[4084-:12]))) & (CSRAdrM != MTIMEH))
				CSRCReadValM = HPMCOUNTERH_REGW[CounterNumM];
			else if (((CSRAdrM >= HPMCOUNTERHBASE) & (CSRAdrM < (HPMCOUNTERHBASE + P[4084-:12]))) & ~CSRWriteM)
				CSRCReadValM = HPMCOUNTERH_REGW[CounterNumM];
			else begin
				CSRCReadValM = 1'sb0;
				IllegalCSRCAccessM = 1'b1;
			end
		end
		else begin
			CSRCReadValM = 1'sb0;
			IllegalCSRCAccessM = 1'b1;
		end
	end
	initial _sv2v_0 = 0;
endmodule
module csri (
	clk,
	reset,
	CSRMWriteM,
	CSRSWriteM,
	CSRWriteValM,
	CSRAdrM,
	MExtInt,
	SExtInt,
	MTimerInt,
	STimerInt,
	MSwInt,
	MIDELEG_REGW,
	ENVCFG_STCE,
	MIP_REGW,
	MIE_REGW,
	MIP_REGW_writeable
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire CSRMWriteM;
	input wire CSRSWriteM;
	input wire [$signed(P[4216-:32]) - 1:0] CSRWriteValM;
	input wire [11:0] CSRAdrM;
	input wire MExtInt;
	input wire SExtInt;
	input wire MTimerInt;
	input wire STimerInt;
	input wire MSwInt;
	input wire [11:0] MIDELEG_REGW;
	input wire ENVCFG_STCE;
	output wire [11:0] MIP_REGW;
	output reg [11:0] MIE_REGW;
	output reg [11:0] MIP_REGW_writeable;
	wire [11:0] MIP_WRITE_MASK;
	wire [11:0] SIP_WRITE_MASK;
	wire [11:0] MIE_WRITE_MASK;
	wire WriteMIPM;
	wire WriteMIEM;
	wire WriteSIPM;
	wire WriteSIEM;
	wire STIP;
	localparam MIE = 12'h304;
	localparam MIP = 12'h344;
	localparam SIE = 12'h104;
	localparam SIP = 12'h144;
	assign WriteMIPM = CSRMWriteM & (CSRAdrM == MIP);
	assign WriteMIEM = CSRMWriteM & (CSRAdrM == MIE);
	assign WriteSIPM = CSRSWriteM & (CSRAdrM == SIP);
	assign WriteSIEM = CSRSWriteM & (CSRAdrM == SIE);
	generate
		if (P[1487]) begin : mask
			if (P[4068]) begin : genblk1
				assign MIP_WRITE_MASK = (ENVCFG_STCE ? 12'h202 : 12'h222);
				assign STIP = (ENVCFG_STCE ? STimerInt : MIP_REGW_writeable[5]);
			end
			else begin : genblk1
				assign MIP_WRITE_MASK = 12'h222;
				assign STIP = MIP_REGW_writeable[5];
			end
			assign SIP_WRITE_MASK = 12'h002 & MIDELEG_REGW;
			assign MIE_WRITE_MASK = 12'haaa;
		end
		else begin : mask
			assign MIP_WRITE_MASK = 12'h000;
			assign SIP_WRITE_MASK = 12'h000;
			assign MIE_WRITE_MASK = 12'h888;
			assign STIP = 1'sb0;
		end
	endgenerate
	always @(posedge clk)
		if (reset)
			MIP_REGW_writeable <= 12'b000000000000;
		else if (WriteMIPM)
			MIP_REGW_writeable <= CSRWriteValM[11:0] & MIP_WRITE_MASK;
		else if (WriteSIPM)
			MIP_REGW_writeable <= (CSRWriteValM[11:0] & SIP_WRITE_MASK) | (MIP_REGW_writeable & ~SIP_WRITE_MASK);
	always @(posedge clk)
		if (reset)
			MIE_REGW <= 12'b000000000000;
		else if (WriteMIEM)
			MIE_REGW <= CSRWriteValM[11:0] & MIE_WRITE_MASK;
		else if (WriteSIEM)
			MIE_REGW <= ((CSRWriteValM[11:0] & 12'h222) & MIDELEG_REGW) | (MIE_REGW & 12'h888);
	assign MIP_REGW = {MExtInt, 1'b0, SExtInt | MIP_REGW_writeable[9], 1'b0, MTimerInt, 1'b0, STIP, 1'b0, MSwInt, 1'b0, MIP_REGW_writeable[1], 1'b0};
endmodule
module csrm (
	clk,
	reset,
	UngatedCSRMWriteM,
	CSRMWriteM,
	MTrapM,
	CSRAdrM,
	NextEPCM,
	NextMtvalM,
	MSTATUS_REGW,
	MSTATUSH_REGW,
	NextCauseM,
	CSRWriteValM,
	MIP_REGW,
	MIE_REGW,
	CSRMReadValM,
	MTVEC_REGW,
	MEPC_REGW,
	MCOUNTEREN_REGW,
	MCOUNTINHIBIT_REGW,
	MEDELEG_REGW,
	MIDELEG_REGW,
	PMPCFG_ARRAY_REGW,
	PMPADDR_ARRAY_REGW,
	WriteMSTATUSM,
	WriteMSTATUSHM,
	IllegalCSRMAccessM,
	IllegalCSRMWriteReadonlyM,
	MENVCFG_REGW
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire UngatedCSRMWriteM;
	input wire CSRMWriteM;
	input wire MTrapM;
	input wire [11:0] CSRAdrM;
	input wire [$signed(P[4216-:32]) - 1:0] NextEPCM;
	input wire [$signed(P[4216-:32]) - 1:0] NextMtvalM;
	input wire [$signed(P[4216-:32]) - 1:0] MSTATUS_REGW;
	input wire [$signed(P[4216-:32]) - 1:0] MSTATUSH_REGW;
	input wire [4:0] NextCauseM;
	input wire [$signed(P[4216-:32]) - 1:0] CSRWriteValM;
	input wire [11:0] MIP_REGW;
	input wire [11:0] MIE_REGW;
	output reg [$signed(P[4216-:32]) - 1:0] CSRMReadValM;
	output wire [$signed(P[4216-:32]) - 1:0] MTVEC_REGW;
	output wire [$signed(P[4216-:32]) - 1:0] MEPC_REGW;
	output wire [31:0] MCOUNTEREN_REGW;
	output wire [31:0] MCOUNTINHIBIT_REGW;
	output wire [15:0] MEDELEG_REGW;
	output wire [11:0] MIDELEG_REGW;
	output wire [($signed(P[3728-:32]) * 8) - 1:0] PMPCFG_ARRAY_REGW;
	output wire [(($signed(P[1640-:32]) - 3) >= 0 ? ($signed(P[3728-:32]) * ($signed(P[1640-:32]) - 2)) - 1 : ($signed(P[3728-:32]) * (4 - $signed(P[1640-:32]))) + ($signed(P[1640-:32]) - 4)):(($signed(P[1640-:32]) - 3) >= 0 ? 0 : $signed(P[1640-:32]) - 3)] PMPADDR_ARRAY_REGW;
	output wire WriteMSTATUSM;
	output wire WriteMSTATUSHM;
	output reg IllegalCSRMAccessM;
	output wire IllegalCSRMWriteReadonlyM;
	output wire [63:0] MENVCFG_REGW;
	wire [$signed(P[4216-:32]) - 1:0] MISA_REGW;
	wire [$signed(P[4216-:32]) - 1:0] MHARTID_REGW;
	wire [$signed(P[4216-:32]) - 1:0] MSCRATCH_REGW;
	wire [$signed(P[4216-:32]) - 1:0] MTVAL_REGW;
	wire [$signed(P[4216-:32]) - 1:0] MCAUSE_REGW;
	wire [$signed(P[4216-:32]) - 1:0] MENVCFGH_REGW;
	wire [$signed(P[4216-:32]) - 1:0] TVECWriteValM;
	wire WriteMTVECM;
	wire WriteMEDELEGM;
	wire WriteMIDELEGM;
	wire WriteMSCRATCHM;
	wire WriteMEPCM;
	wire WriteMCAUSEM;
	wire WriteMTVALM;
	wire WriteMCOUNTERENM;
	wire WriteMCOUNTINHIBITM;
	localparam MVENDORID = 12'hf11;
	localparam MARCHID = 12'hf12;
	localparam MIMPID = 12'hf13;
	localparam MHARTID = 12'hf14;
	localparam MCONFIGPTR = 12'hf15;
	localparam MSTATUS = 12'h300;
	localparam MISA_ADR = 12'h301;
	localparam MEDELEG = 12'h302;
	localparam MIDELEG = 12'h303;
	localparam MIE = 12'h304;
	localparam MTVEC = 12'h305;
	localparam MCOUNTEREN = 12'h306;
	localparam MENVCFG = 12'h30a;
	localparam MSTATUSH = 12'h310;
	localparam MENVCFGH = 12'h31a;
	localparam MCOUNTINHIBIT = 12'h320;
	localparam MSCRATCH = 12'h340;
	localparam MEPC = 12'h341;
	localparam MCAUSE = 12'h342;
	localparam MTVAL = 12'h343;
	localparam MIP = 12'h344;
	localparam PMPCFG0 = 12'h3a0;
	localparam PMPADDR0 = 12'h3b0;
	localparam TSELECT = 12'h7a0;
	localparam TDATA1 = 12'h7a1;
	localparam TDATA2 = 12'h7a2;
	localparam TDATA3 = 12'h7a3;
	localparam DCSR = 12'h7b0;
	localparam DPC = 12'h7b1;
	localparam DSCRATCH0 = 12'h7b2;
	localparam DSCRATCH1 = 12'h7b3;
	localparam ZERO = {$signed(P[4216-:32]) {1'b0}};
	localparam MEDELEG_MASK = (P[1754] ? 16'hb3fe : 16'hb3ff);
	localparam MIDELEG_MASK = 12'h222;
	genvar _gv_i_5;
	generate
		if ($signed(P[3728-:32]) > 0) begin : pmp
			wire [$signed(P[3728-:32]) - 1:0] WritePMPCFGM;
			wire [$signed(P[3728-:32]) - 1:0] WritePMPADDRM;
			wire [7:0] CSRPMPWriteValM [$signed(P[3728-:32]) - 1:0];
			wire [7:0] CSRPMPLegalizedWriteValM [$signed(P[3728-:32]) - 1:0];
			wire [1:0] CSRPMPWRLegalizedWriteValM [$signed(P[3728-:32]) - 1:0];
			wire [$signed(P[3728-:32]) - 1:0] ADDRLocked;
			wire [$signed(P[3728-:32]) - 1:0] CFGLocked;
			for (_gv_i_5 = 0; _gv_i_5 < $signed(P[3728-:32]); _gv_i_5 = _gv_i_5 + 1) begin : genblk1
				localparam i = _gv_i_5;
				assign CFGLocked[i] = PMPCFG_ARRAY_REGW[(i * 8) + 7];
				if (i == ($signed(P[3728-:32]) - 1)) begin : genblk1
					assign ADDRLocked[i] = PMPCFG_ARRAY_REGW[(i * 8) + 7];
				end
				else begin : genblk1
					assign ADDRLocked[i] = PMPCFG_ARRAY_REGW[(i * 8) + 7] | (PMPCFG_ARRAY_REGW[((i + 1) * 8) + 7] & (PMPCFG_ARRAY_REGW[((i + 1) * 8) + 4-:2] == 2'b01));
				end
				assign WritePMPADDRM[i] = (CSRMWriteM & (CSRAdrM == (PMPADDR0 + i))) & ~ADDRLocked[i];
				flopenr #(.WIDTH($signed(P[1640-:32]) - 2)) PMPADDRreg(
					.clk(clk),
					.reset(reset),
					.en(WritePMPADDRM[i]),
					.d(CSRWriteValM[$signed(P[1640-:32]) - 3:0]),
					.q(PMPADDR_ARRAY_REGW[(($signed(P[1640-:32]) - 3) >= 0 ? 0 : $signed(P[1640-:32]) - 3) + (i * (($signed(P[1640-:32]) - 3) >= 0 ? $signed(P[1640-:32]) - 2 : 4 - $signed(P[1640-:32])))+:(($signed(P[1640-:32]) - 3) >= 0 ? $signed(P[1640-:32]) - 2 : 4 - $signed(P[1640-:32]))])
				);
				if ($signed(P[4216-:32]) == 64) begin : genblk2
					assign WritePMPCFGM[i] = (CSRMWriteM & (CSRAdrM == (PMPCFG0 + (2 * (i / 8))))) & ~CFGLocked[i];
					assign CSRPMPWriteValM[i] = CSRWriteValM[((i % 8) * 8) + 7:(i % 8) * 8];
				end
				else begin : genblk2
					assign WritePMPCFGM[i] = (CSRMWriteM & (CSRAdrM == (PMPCFG0 + (i / 4)))) & ~CFGLocked[i];
					assign CSRPMPWriteValM[i] = CSRWriteValM[((i % 4) * 8) + 7:(i % 4) * 8];
				end
				assign CSRPMPWRLegalizedWriteValM[i] = {CSRPMPWriteValM[i][1] & CSRPMPWriteValM[i][0], CSRPMPWriteValM[i][0]};
				assign CSRPMPLegalizedWriteValM[i] = {CSRPMPWriteValM[i][7], 2'b00, CSRPMPWriteValM[i][4:2], CSRPMPWRLegalizedWriteValM[i]};
				flopenr #(.WIDTH(8)) PMPCFGreg(
					.clk(clk),
					.reset(reset),
					.en(WritePMPCFGM[i]),
					.d(CSRPMPLegalizedWriteValM[i]),
					.q(PMPCFG_ARRAY_REGW[i * 8+:8])
				);
			end
		end
	endgenerate
	localparam MISA_26 = $unsigned($signed(P[4183-:32])) & 32'h03ffffff;
	assign MISA_REGW = {($signed(P[4216-:32]) == 32 ? 2'b01 : 2'b10), {$signed(P[4216-:32]) - 28 {1'b0}}, MISA_26[25:0]};
	assign MHARTID_REGW = 1'sb0;
	assign WriteMSTATUSM = CSRMWriteM & (CSRAdrM == MSTATUS);
	assign WriteMSTATUSHM = (CSRMWriteM & (CSRAdrM == MSTATUSH)) & ($signed(P[4216-:32]) == 32);
	assign WriteMTVECM = CSRMWriteM & (CSRAdrM == MTVEC);
	assign WriteMEDELEGM = CSRMWriteM & (CSRAdrM == MEDELEG);
	assign WriteMIDELEGM = CSRMWriteM & (CSRAdrM == MIDELEG);
	assign WriteMSCRATCHM = CSRMWriteM & (CSRAdrM == MSCRATCH);
	assign WriteMEPCM = MTrapM | (CSRMWriteM & (CSRAdrM == MEPC));
	assign WriteMCAUSEM = MTrapM | (CSRMWriteM & (CSRAdrM == MCAUSE));
	assign WriteMTVALM = MTrapM | (CSRMWriteM & (CSRAdrM == MTVAL));
	assign WriteMCOUNTERENM = CSRMWriteM & (CSRAdrM == MCOUNTEREN);
	assign WriteMCOUNTINHIBITM = CSRMWriteM & (CSRAdrM == MCOUNTINHIBIT);
	assign IllegalCSRMWriteReadonlyM = UngatedCSRMWriteM & (((((CSRAdrM == MVENDORID) | (CSRAdrM == MARCHID)) | (CSRAdrM == MIMPID)) | (CSRAdrM == MHARTID)) | (CSRAdrM == MCONFIGPTR));
	assign TVECWriteValM = (CSRWriteValM[0] ? {CSRWriteValM[$signed(P[4216-:32]) - 1:6], 6'b000001} : {CSRWriteValM[$signed(P[4216-:32]) - 1:2], 2'b00});
	flopenr #(.WIDTH($signed(P[4216-:32]))) MTVECreg(
		.clk(clk),
		.reset(reset),
		.en(WriteMTVECM),
		.d(TVECWriteValM),
		.q(MTVEC_REGW)
	);
	generate
		if (P[1487]) begin : deleg
			flopenr #(.WIDTH(16)) MEDELEGreg(
				.clk(clk),
				.reset(reset),
				.en(WriteMEDELEGM),
				.d(CSRWriteValM[15:0] & MEDELEG_MASK),
				.q(MEDELEG_REGW)
			);
			flopenr #(.WIDTH(12)) MIDELEGreg(
				.clk(clk),
				.reset(reset),
				.en(WriteMIDELEGM),
				.d(CSRWriteValM[11:0] & MIDELEG_MASK),
				.q(MIDELEG_REGW)
			);
		end
		else begin : genblk2
			assign {MEDELEG_REGW, MIDELEG_REGW} = 1'sb0;
		end
	endgenerate
	flopenr #(.WIDTH($signed(P[4216-:32]))) MSCRATCHreg(
		.clk(clk),
		.reset(reset),
		.en(WriteMSCRATCHM),
		.d(CSRWriteValM),
		.q(MSCRATCH_REGW)
	);
	flopenr #(.WIDTH($signed(P[4216-:32]))) MEPCreg(
		.clk(clk),
		.reset(reset),
		.en(WriteMEPCM),
		.d(NextEPCM),
		.q(MEPC_REGW)
	);
	flopenr #(.WIDTH($signed(P[4216-:32]))) MCAUSEreg(
		.clk(clk),
		.reset(reset),
		.en(WriteMCAUSEM),
		.d({NextCauseM[4], {$signed(P[4216-:32]) - 5 {1'b0}}, NextCauseM[3:0]}),
		.q(MCAUSE_REGW)
	);
	flopenr #(.WIDTH($signed(P[4216-:32]))) MTVALreg(
		.clk(clk),
		.reset(reset),
		.en(WriteMTVALM),
		.d(NextMtvalM),
		.q(MTVAL_REGW)
	);
	flopenr #(.WIDTH(32)) MCOUNTINHIBITreg(
		.clk(clk),
		.reset(reset),
		.en(WriteMCOUNTINHIBITM),
		.d({CSRWriteValM[31:2], 1'b0, CSRWriteValM[0]}),
		.q(MCOUNTINHIBIT_REGW)
	);
	generate
		if (P[1486]) begin : mcounteren
			flopenr #(.WIDTH(32)) MCOUNTERENreg(
				.clk(clk),
				.reset(reset),
				.en(WriteMCOUNTERENM),
				.d(CSRWriteValM[31:0]),
				.q(MCOUNTEREN_REGW)
			);
		end
		else begin : genblk3
			assign MCOUNTEREN_REGW = 1'sb0;
		end
		if (P[1486]) begin : genblk4
			wire WriteMENVCFGM;
			wire [63:0] MENVCFG_PreWriteValM;
			wire [63:0] MENVCFG_WriteValM;
			wire [1:0] LegalizedCBIE;
			assign WriteMENVCFGM = CSRMWriteM & (CSRAdrM == MENVCFG);
			assign LegalizedCBIE = (MENVCFG_PreWriteValM[5:4] == 2'b10 ? MENVCFG_REGW[5:4] : MENVCFG_PreWriteValM[5:4]);
			assign MENVCFG_WriteValM = {MENVCFG_PreWriteValM[63] & P[4068], MENVCFG_PreWriteValM[62] & P[4057], MENVCFG_PreWriteValM[61] & P[4064], 53'b00000000000000000000000000000000000000000000000000000, MENVCFG_PreWriteValM[7] & P[4061], MENVCFG_PreWriteValM[6] & P[4062], LegalizedCBIE & {2 {P[4062]}}, 3'b000, (MENVCFG_PreWriteValM[0] & P[1487]) & P[4067]};
			if ($signed(P[4216-:32]) == 64) begin : genblk1
				assign MENVCFG_PreWriteValM = CSRWriteValM;
				flopenr #(.WIDTH($signed(P[4216-:32]))) MENVCFGreg(
					.clk(clk),
					.reset(reset),
					.en(WriteMENVCFGM),
					.d(MENVCFG_WriteValM),
					.q(MENVCFG_REGW)
				);
				assign MENVCFGH_REGW = 1'sb0;
			end
			else begin : genblk1
				wire WriteMENVCFGHM;
				assign MENVCFG_PreWriteValM = {CSRWriteValM, CSRWriteValM};
				assign WriteMENVCFGHM = (CSRMWriteM & (CSRAdrM == MENVCFGH)) & ($signed(P[4216-:32]) == 32);
				flopenr #(.WIDTH($signed(P[4216-:32]))) MENVCFGreg(
					.clk(clk),
					.reset(reset),
					.en(WriteMENVCFGM),
					.d(MENVCFG_WriteValM[31:0]),
					.q(MENVCFG_REGW[31:0])
				);
				flopenr #(.WIDTH($signed(P[4216-:32]))) MENVCFGHreg(
					.clk(clk),
					.reset(reset),
					.en(WriteMENVCFGHM),
					.d(MENVCFG_WriteValM[63:32]),
					.q(MENVCFG_REGW[63:32])
				);
				assign MENVCFGH_REGW = MENVCFG_REGW[63:32];
			end
		end
		else begin : genblk4
			assign MENVCFG_REGW = 1'sb0;
			assign MENVCFGH_REGW = 1'sb0;
		end
	endgenerate
	reg [5:0] entry;
	always @(*) begin
		if (_sv2v_0)
			;
		entry = 1'sb0;
		CSRMReadValM = 1'sb0;
		IllegalCSRMAccessM = !P[1487] & ((CSRAdrM == MEDELEG) | (CSRAdrM == MIDELEG));
		if (($unsigned(CSRAdrM) >= PMPADDR0) & ($unsigned(CSRAdrM) < (PMPADDR0 + $signed(P[3728-:32]))))
			CSRMReadValM = {{$signed(P[4216-:32]) - ($signed(P[1640-:32]) - 2) {1'b0}}, PMPADDR_ARRAY_REGW[(($signed(P[1640-:32]) - 3) >= 0 ? 0 : $signed(P[1640-:32]) - 3) + ((CSRAdrM - PMPADDR0) * (($signed(P[1640-:32]) - 3) >= 0 ? $signed(P[1640-:32]) - 2 : 4 - $signed(P[1640-:32])))+:(($signed(P[1640-:32]) - 3) >= 0 ? $signed(P[1640-:32]) - 2 : 4 - $signed(P[1640-:32]))]};
		else if ((($unsigned(CSRAdrM) >= PMPCFG0) & ($unsigned(CSRAdrM) < (PMPCFG0 + ($signed(P[3728-:32]) / 4)))) & (($signed(P[4216-:32]) == 32) | (CSRAdrM[0] == 0))) begin
			if ($signed(P[4216-:32]) == 64) begin
				entry = ({CSRAdrM[11:1], 1'b0} - PMPCFG0) * 4;
				CSRMReadValM = {PMPCFG_ARRAY_REGW[(entry + 7) * 8+:8], PMPCFG_ARRAY_REGW[(entry + 6) * 8+:8], PMPCFG_ARRAY_REGW[(entry + 5) * 8+:8], PMPCFG_ARRAY_REGW[(entry + 4) * 8+:8], PMPCFG_ARRAY_REGW[(entry + 3) * 8+:8], PMPCFG_ARRAY_REGW[(entry + 2) * 8+:8], PMPCFG_ARRAY_REGW[(entry + 1) * 8+:8], PMPCFG_ARRAY_REGW[entry * 8+:8]};
			end
			else begin
				entry = (CSRAdrM - PMPCFG0) * 4;
				CSRMReadValM = {PMPCFG_ARRAY_REGW[(entry + 3) * 8+:8], PMPCFG_ARRAY_REGW[(entry + 2) * 8+:8], PMPCFG_ARRAY_REGW[(entry + 1) * 8+:8], PMPCFG_ARRAY_REGW[entry * 8+:8]};
			end
		end
		else
			case (CSRAdrM)
				MISA_ADR: CSRMReadValM = MISA_REGW;
				MVENDORID: CSRMReadValM = {{$signed(P[4216-:32]) - 32 {1'b0}}, 32'h00000602};
				MARCHID: CSRMReadValM = {{$signed(P[4216-:32]) - 32 {1'b0}}, 32'h00000024};
				MIMPID: CSRMReadValM = {{$signed(P[4216-:32]) - 12 {1'b0}}, 12'h100};
				MHARTID: CSRMReadValM = MHARTID_REGW;
				MCONFIGPTR: CSRMReadValM = 1'sb0;
				MSTATUS: CSRMReadValM = MSTATUS_REGW;
				MSTATUSH:
					if ($signed(P[4216-:32]) == 32)
						CSRMReadValM = MSTATUSH_REGW;
					else
						IllegalCSRMAccessM = 1'b1;
				MTVEC: CSRMReadValM = MTVEC_REGW;
				MEDELEG: CSRMReadValM = {{$signed(P[4216-:32]) - 16 {1'b0}}, MEDELEG_REGW};
				MIDELEG: CSRMReadValM = {{$signed(P[4216-:32]) - 12 {1'b0}}, MIDELEG_REGW};
				MIP: CSRMReadValM = {{$signed(P[4216-:32]) - 12 {1'b0}}, MIP_REGW};
				MIE: CSRMReadValM = {{$signed(P[4216-:32]) - 12 {1'b0}}, MIE_REGW};
				MSCRATCH: CSRMReadValM = MSCRATCH_REGW;
				MEPC: CSRMReadValM = MEPC_REGW;
				MCAUSE: CSRMReadValM = MCAUSE_REGW;
				MTVAL: CSRMReadValM = MTVAL_REGW;
				MCOUNTEREN: CSRMReadValM = {{$signed(P[4216-:32]) - 32 {1'b0}}, MCOUNTEREN_REGW};
				MENVCFG:
					if (P[1486])
						CSRMReadValM = MENVCFG_REGW[$signed(P[4216-:32]) - 1:0];
					else
						IllegalCSRMAccessM = 1'b1;
				MENVCFGH:
					if (P[1486] & ($signed(P[4216-:32]) == 32))
						CSRMReadValM = MENVCFGH_REGW;
					else
						IllegalCSRMAccessM = 1'b1;
				MCOUNTINHIBIT: CSRMReadValM = {{$signed(P[4216-:32]) - 32 {1'b0}}, MCOUNTINHIBIT_REGW};
				default: IllegalCSRMAccessM = 1'b1;
			endcase
	end
	initial _sv2v_0 = 0;
endmodule
module csrs (
	clk,
	reset,
	CSRSWriteM,
	STrapM,
	CSRAdrM,
	NextEPCM,
	NextMtvalM,
	SSTATUS_REGW,
	NextCauseM,
	STATUS_TVM,
	CSRWriteValM,
	PrivilegeModeW,
	CSRSReadValM,
	STVEC_REGW,
	SEPC_REGW,
	SCOUNTEREN_REGW,
	SATP_REGW,
	MIP_REGW,
	MIE_REGW,
	MIDELEG_REGW,
	MTIME_CLINT,
	STCE,
	WriteSSTATUSM,
	IllegalCSRSAccessM,
	STimerInt,
	SENVCFG_REGW
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire CSRSWriteM;
	input wire STrapM;
	input wire [11:0] CSRAdrM;
	input wire [$signed(P[4216-:32]) - 1:0] NextEPCM;
	input wire [$signed(P[4216-:32]) - 1:0] NextMtvalM;
	input wire [$signed(P[4216-:32]) - 1:0] SSTATUS_REGW;
	input wire [4:0] NextCauseM;
	input wire STATUS_TVM;
	input wire [$signed(P[4216-:32]) - 1:0] CSRWriteValM;
	input wire [1:0] PrivilegeModeW;
	output reg [$signed(P[4216-:32]) - 1:0] CSRSReadValM;
	output wire [$signed(P[4216-:32]) - 1:0] STVEC_REGW;
	output wire [$signed(P[4216-:32]) - 1:0] SEPC_REGW;
	output wire [31:0] SCOUNTEREN_REGW;
	output wire [$signed(P[4216-:32]) - 1:0] SATP_REGW;
	input wire [11:0] MIP_REGW;
	input wire [11:0] MIE_REGW;
	input wire [11:0] MIDELEG_REGW;
	input wire [63:0] MTIME_CLINT;
	input wire STCE;
	output wire WriteSSTATUSM;
	output reg IllegalCSRSAccessM;
	output wire STimerInt;
	output wire [$signed(P[4216-:32]) - 1:0] SENVCFG_REGW;
	localparam SSTATUS = 12'h100;
	localparam SIE = 12'h104;
	localparam STVEC = 12'h105;
	localparam SCOUNTEREN = 12'h106;
	localparam SENVCFG = 12'h10a;
	localparam SSCRATCH = 12'h140;
	localparam SEPC = 12'h141;
	localparam SCAUSE = 12'h142;
	localparam STVAL = 12'h143;
	localparam SIP = 12'h144;
	localparam STIMECMP = 12'h14d;
	localparam STIMECMPH = 12'h15d;
	localparam SATP = 12'h180;
	wire WriteSTVECM;
	wire WriteSSCRATCHM;
	wire WriteSEPCM;
	wire WriteSCAUSEM;
	wire WriteSTVALM;
	wire WriteSATPM;
	wire WriteSCOUNTERENM;
	wire WriteSTIMECMPM;
	wire WriteSTIMECMPHM;
	wire WriteSENVCFGM;
	wire [$signed(P[4216-:32]) - 1:0] SSCRATCH_REGW;
	wire [$signed(P[4216-:32]) - 1:0] STVAL_REGW;
	wire [$signed(P[4216-:32]) - 1:0] SCAUSE_REGW;
	wire [$signed(P[4216-:32]) - 1:0] SENVCFG_WriteValM;
	wire [$signed(P[4216-:32]) - 1:0] TVECWriteValM;
	wire [63:0] STIMECMP_REGW;
	assign WriteSSTATUSM = CSRSWriteM & (CSRAdrM == SSTATUS);
	assign WriteSTVECM = CSRSWriteM & (CSRAdrM == STVEC);
	assign WriteSSCRATCHM = CSRSWriteM & (CSRAdrM == SSCRATCH);
	assign WriteSEPCM = STrapM | (CSRSWriteM & (CSRAdrM == SEPC));
	assign WriteSCAUSEM = STrapM | (CSRSWriteM & (CSRAdrM == SCAUSE));
	assign WriteSTVALM = STrapM | (CSRSWriteM & (CSRAdrM == STVAL));
	generate
		if ($signed(P[4216-:32]) == 64) begin : genblk1
			wire LegalSatpModeM;
			assign LegalSatpModeM = P[4067] & (((CSRWriteValM[63:60] == 0) | (CSRWriteValM[63:60] == P[1504-:4])) | (CSRWriteValM[63:60] == P[1500-:4]));
			assign WriteSATPM = ((CSRSWriteM & (CSRAdrM == SATP)) & ((PrivilegeModeW == P[1742-:2]) | ~STATUS_TVM)) & LegalSatpModeM;
		end
		else begin : genblk1
			assign WriteSATPM = ((CSRSWriteM & (CSRAdrM == SATP)) & ((PrivilegeModeW == P[1742-:2]) | ~STATUS_TVM)) & P[4067];
		end
	endgenerate
	assign WriteSCOUNTERENM = CSRSWriteM & (CSRAdrM == SCOUNTEREN);
	assign WriteSENVCFGM = CSRSWriteM & (CSRAdrM == SENVCFG);
	assign WriteSTIMECMPM = (CSRSWriteM & (CSRAdrM == STIMECMP)) & STCE;
	assign WriteSTIMECMPHM = ((CSRSWriteM & (CSRAdrM == STIMECMPH)) & STCE) & ($signed(P[4216-:32]) == 32);
	assign TVECWriteValM = (CSRWriteValM[0] ? {CSRWriteValM[$signed(P[4216-:32]) - 1:6], 6'b000001} : {CSRWriteValM[$signed(P[4216-:32]) - 1:2], 2'b00});
	flopenr #(.WIDTH($signed(P[4216-:32]))) STVECreg(
		.clk(clk),
		.reset(reset),
		.en(WriteSTVECM),
		.d(TVECWriteValM),
		.q(STVEC_REGW)
	);
	flopenr #(.WIDTH($signed(P[4216-:32]))) SSCRATCHreg(
		.clk(clk),
		.reset(reset),
		.en(WriteSSCRATCHM),
		.d(CSRWriteValM),
		.q(SSCRATCH_REGW)
	);
	flopenr #(.WIDTH($signed(P[4216-:32]))) SEPCreg(
		.clk(clk),
		.reset(reset),
		.en(WriteSEPCM),
		.d(NextEPCM),
		.q(SEPC_REGW)
	);
	flopenr #(.WIDTH($signed(P[4216-:32]))) SCAUSEreg(
		.clk(clk),
		.reset(reset),
		.en(WriteSCAUSEM),
		.d({NextCauseM[4], {$signed(P[4216-:32]) - 5 {1'b0}}, NextCauseM[3:0]}),
		.q(SCAUSE_REGW)
	);
	flopenr #(.WIDTH($signed(P[4216-:32]))) STVALreg(
		.clk(clk),
		.reset(reset),
		.en(WriteSTVALM),
		.d(NextMtvalM),
		.q(STVAL_REGW)
	);
	generate
		if (P[4067]) begin : genblk2
			flopenr #(.WIDTH($signed(P[4216-:32]))) SATPreg(
				.clk(clk),
				.reset(reset),
				.en(WriteSATPM),
				.d(CSRWriteValM),
				.q(SATP_REGW)
			);
		end
		else begin : genblk2
			assign SATP_REGW = 1'sb0;
		end
	endgenerate
	flopenr #(.WIDTH(32)) SCOUNTERENreg(
		.clk(clk),
		.reset(reset),
		.en(WriteSCOUNTERENM),
		.d(CSRWriteValM[31:0]),
		.q(SCOUNTEREN_REGW)
	);
	generate
		if (P[4068]) begin : sstc
			if ($signed(P[4216-:32]) == 64) begin : sstc64
				flopenr #(.WIDTH($signed(P[4216-:32]))) STIMECMPreg(
					.clk(clk),
					.reset(reset),
					.en(WriteSTIMECMPM),
					.d(CSRWriteValM),
					.q(STIMECMP_REGW)
				);
			end
			else begin : sstc32
				flopenr #(.WIDTH($signed(P[4216-:32]))) STIMECMPreg(
					.clk(clk),
					.reset(reset),
					.en(WriteSTIMECMPM),
					.d(CSRWriteValM),
					.q(STIMECMP_REGW[31:0])
				);
				flopenr #(.WIDTH($signed(P[4216-:32]))) STIMECMPHreg(
					.clk(clk),
					.reset(reset),
					.en(WriteSTIMECMPHM),
					.d(CSRWriteValM),
					.q(STIMECMP_REGW[63:32])
				);
			end
		end
		else begin : genblk3
			assign STIMECMP_REGW = 1'sb0;
		end
		if (P[4068]) begin : genblk4
			assign STimerInt = {1'b0, MTIME_CLINT} >= {1'b0, STIMECMP_REGW};
		end
		else begin : genblk4
			assign STimerInt = 1'b0;
		end
	endgenerate
	wire [1:0] LegalizedCBIE;
	assign LegalizedCBIE = (CSRWriteValM[5:4] == 2'b10 ? SENVCFG_REGW[5:4] : CSRWriteValM[5:4]);
	assign SENVCFG_WriteValM = {{$signed(P[4216-:32]) - 8 {1'b0}}, CSRWriteValM[7] & P[4061], CSRWriteValM[6] & P[4062], LegalizedCBIE & {2 {P[4062]}}, 3'b000, CSRWriteValM[0] & P[4067]};
	flopenr #(.WIDTH($signed(P[4216-:32]))) SENVCFGreg(
		.clk(clk),
		.reset(reset),
		.en(WriteSENVCFGM),
		.d(SENVCFG_WriteValM),
		.q(SENVCFG_REGW)
	);
	always @(*) begin : csrr
		if (_sv2v_0)
			;
		IllegalCSRSAccessM = 1'b0;
		case (CSRAdrM)
			SSTATUS: CSRSReadValM = SSTATUS_REGW;
			STVEC: CSRSReadValM = STVEC_REGW;
			SIP: CSRSReadValM = {{$signed(P[4216-:32]) - 12 {1'b0}}, (MIP_REGW & 12'h222) & MIDELEG_REGW};
			SIE: CSRSReadValM = {{$signed(P[4216-:32]) - 12 {1'b0}}, (MIE_REGW & 12'h222) & MIDELEG_REGW};
			SSCRATCH: CSRSReadValM = SSCRATCH_REGW;
			SEPC: CSRSReadValM = SEPC_REGW;
			SCAUSE: CSRSReadValM = SCAUSE_REGW;
			STVAL: CSRSReadValM = STVAL_REGW;
			SATP:
				if (P[4067] & ((PrivilegeModeW == P[1742-:2]) | ~STATUS_TVM))
					CSRSReadValM = SATP_REGW;
				else begin
					CSRSReadValM = 1'sb0;
					IllegalCSRSAccessM = 1'b1;
				end
			SCOUNTEREN: CSRSReadValM = {{$signed(P[4216-:32]) - 32 {1'b0}}, SCOUNTEREN_REGW};
			SENVCFG: CSRSReadValM = SENVCFG_REGW;
			STIMECMP:
				if (STCE)
					CSRSReadValM = STIMECMP_REGW[$signed(P[4216-:32]) - 1:0];
				else begin
					CSRSReadValM = 1'sb0;
					IllegalCSRSAccessM = 1'b1;
				end
			STIMECMPH:
				if (STCE & ($signed(P[4216-:32]) == 32))
					CSRSReadValM = {{$signed(P[4216-:32]) - 32 {1'b0}}, STIMECMP_REGW[63:32]};
				else begin
					CSRSReadValM = 1'sb0;
					IllegalCSRSAccessM = 1'b1;
				end
			default: begin
				CSRSReadValM = 1'sb0;
				IllegalCSRSAccessM = 1'b1;
			end
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
module csrsr (
	clk,
	reset,
	StallW,
	WriteMSTATUSM,
	WriteMSTATUSHM,
	WriteSSTATUSM,
	TrapM,
	FRegWriteM,
	NextPrivilegeModeM,
	PrivilegeModeW,
	mretM,
	sretM,
	WriteFRMM,
	SetOrWriteFFLAGSM,
	CSRWriteValM,
	SelHPTW,
	MSTATUS_REGW,
	SSTATUS_REGW,
	MSTATUSH_REGW,
	STATUS_MPP,
	STATUS_SPP,
	STATUS_TSR,
	STATUS_TW,
	STATUS_MIE,
	STATUS_SIE,
	STATUS_MXR,
	STATUS_SUM,
	STATUS_MPRV,
	STATUS_TVM,
	STATUS_FS,
	BigEndianM
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallW;
	input wire WriteMSTATUSM;
	input wire WriteMSTATUSHM;
	input wire WriteSSTATUSM;
	input wire TrapM;
	input wire FRegWriteM;
	input wire [1:0] NextPrivilegeModeM;
	input wire [1:0] PrivilegeModeW;
	input wire mretM;
	input wire sretM;
	input wire WriteFRMM;
	input wire SetOrWriteFFLAGSM;
	input wire [$signed(P[4216-:32]) - 1:0] CSRWriteValM;
	input wire SelHPTW;
	output wire [$signed(P[4216-:32]) - 1:0] MSTATUS_REGW;
	output wire [$signed(P[4216-:32]) - 1:0] SSTATUS_REGW;
	output wire [$signed(P[4216-:32]) - 1:0] MSTATUSH_REGW;
	output reg [1:0] STATUS_MPP;
	output reg STATUS_SPP;
	output wire STATUS_TSR;
	output wire STATUS_TW;
	output reg STATUS_MIE;
	output reg STATUS_SIE;
	output wire STATUS_MXR;
	output wire STATUS_SUM;
	output wire STATUS_MPRV;
	output wire STATUS_TVM;
	output wire [1:0] STATUS_FS;
	output reg BigEndianM;
	wire STATUS_SD;
	reg STATUS_TW_INT;
	reg STATUS_TSR_INT;
	reg STATUS_TVM_INT;
	reg STATUS_MXR_INT;
	reg STATUS_SUM_INT;
	reg STATUS_MPRV_INT;
	wire [1:0] STATUS_SXL;
	wire [1:0] STATUS_UXL;
	wire [1:0] STATUS_XS;
	reg [1:0] STATUS_FS_INT;
	reg [1:0] STATUS_MPP_NEXT;
	reg STATUS_MPIE;
	reg STATUS_SPIE;
	reg STATUS_UBE;
	reg STATUS_SBE;
	reg STATUS_MBE;
	wire nextMBE;
	wire nextSBE;
	generate
		if ($signed(P[4216-:32]) == 64) begin : csrsr64
			assign MSTATUS_REGW = {STATUS_SD, 25'b0000000000000000000000000, STATUS_MBE, STATUS_SBE, STATUS_SXL, STATUS_UXL, 9'b000000000, STATUS_TSR, STATUS_TW, STATUS_TVM, STATUS_MXR, STATUS_SUM, STATUS_MPRV, STATUS_XS, STATUS_FS, STATUS_MPP, 2'b00, STATUS_SPP, STATUS_MPIE, STATUS_UBE, STATUS_SPIE, 1'b0, STATUS_MIE, 1'b0, STATUS_SIE, 1'b0};
			assign SSTATUS_REGW = {STATUS_SD, 29'b00000000000000000000000000000, STATUS_UXL, 12'b000000000000, STATUS_MXR, STATUS_SUM, 1'b0, STATUS_XS, STATUS_FS, 4'b0000, STATUS_SPP, 1'b0, STATUS_UBE, STATUS_SPIE, 3'b000, STATUS_SIE, 1'b0};
			assign MSTATUSH_REGW = 1'sb0;
		end
		else begin : csrsr32
			assign MSTATUS_REGW = {STATUS_SD, 8'b00000000, STATUS_TSR, STATUS_TW, STATUS_TVM, STATUS_MXR, STATUS_SUM, STATUS_MPRV, STATUS_XS, STATUS_FS, STATUS_MPP, 2'b00, STATUS_SPP, STATUS_MPIE, STATUS_UBE, STATUS_SPIE, 1'b0, STATUS_MIE, 1'b0, STATUS_SIE, 1'b0};
			assign MSTATUSH_REGW = {26'b00000000000000000000000000, STATUS_MBE, STATUS_SBE, 4'b0000};
			assign SSTATUS_REGW = {STATUS_SD, 11'b00000000000, STATUS_MXR, STATUS_SUM, 1'b0, STATUS_XS, STATUS_FS, 4'b0000, STATUS_SPP, 1'b0, STATUS_UBE, STATUS_SPIE, 3'b000, STATUS_SIE, 1'b0};
		end
		if ($signed(P[4216-:32]) == 64) begin : upperstatus
			assign nextMBE = P[4065] & CSRWriteValM[37];
			assign nextSBE = (P[1487] & P[4065]) & CSRWriteValM[36];
		end
		else begin : upperstatus
			assign nextMBE = P[4065] & STATUS_MBE;
			assign nextSBE = (P[1487] & P[4065]) & STATUS_SBE;
		end
	endgenerate
	assign STATUS_TSR = P[1487] & STATUS_TSR_INT;
	assign STATUS_TW = P[1486] & STATUS_TW_INT;
	assign STATUS_TVM = P[1487] & STATUS_TVM_INT;
	assign STATUS_MXR = P[1487] & STATUS_MXR_INT;
	assign STATUS_SXL = (P[1487] ? 2'b10 : 2'b00);
	assign STATUS_UXL = (P[1486] ? 2'b10 : 2'b00);
	assign STATUS_SUM = (P[1487] & P[4067]) & STATUS_SUM_INT;
	assign STATUS_MPRV = P[1486] & STATUS_MPRV_INT;
	assign STATUS_FS = (P[1491] ? STATUS_FS_INT : 2'b00);
	assign STATUS_SD = (STATUS_FS == 2'b11) | (STATUS_XS == 2'b11);
	assign STATUS_XS = 2'b00;
	always @(*) begin
		if (_sv2v_0)
			;
		if ((CSRWriteValM[12:11] == P[1738-:2]) & P[1486])
			STATUS_MPP_NEXT = P[1738-:2];
		else if ((CSRWriteValM[12:11] == P[1740-:2]) & P[1487])
			STATUS_MPP_NEXT = P[1740-:2];
		else if (CSRWriteValM[12:11] == P[1742-:2])
			STATUS_MPP_NEXT = P[1742-:2];
		else
			STATUS_MPP_NEXT = STATUS_MPP;
	end
	generate
		if (P[4065]) begin : endianmux
			reg [1:0] EndiannessPrivMode;
			always @(*) begin
				if (_sv2v_0)
					;
				if (SelHPTW)
					EndiannessPrivMode = P[1740-:2];
				else if ((PrivilegeModeW == P[1742-:2]) & STATUS_MPRV)
					EndiannessPrivMode = STATUS_MPP;
				else
					EndiannessPrivMode = PrivilegeModeW;
				case (EndiannessPrivMode)
					P[1742-:2]: BigEndianM = STATUS_MBE;
					P[1740-:2]: BigEndianM = STATUS_SBE;
					default: BigEndianM = STATUS_UBE;
				endcase
			end
		end
		else begin : endianmux
			wire [1:1] sv2v_tmp_2A6F5;
			assign sv2v_tmp_2A6F5 = 1'b0;
			always @(*) BigEndianM = sv2v_tmp_2A6F5;
		end
	endgenerate
	always @(posedge clk)
		if (reset) begin
			STATUS_TSR_INT <= 1'b0;
			STATUS_TW_INT <= 1'b0;
			STATUS_TVM_INT <= 1'b0;
			STATUS_MXR_INT <= 1'b0;
			STATUS_SUM_INT <= 1'b0;
			STATUS_MPRV_INT <= 1'b0;
			STATUS_FS_INT <= 2'b00;
			STATUS_MPP <= 2'b00;
			STATUS_SPP <= 1'b0;
			STATUS_MPIE <= 1'b0;
			STATUS_SPIE <= 1'b0;
			STATUS_MIE <= 1'b0;
			STATUS_SIE <= 1'b0;
			STATUS_MBE <= 1'b0;
			STATUS_SBE <= 1'b0;
			STATUS_UBE <= 1'b0;
		end
		else if (~StallW) begin
			if (TrapM) begin
				if (NextPrivilegeModeM == P[1742-:2]) begin
					STATUS_MPIE <= STATUS_MIE;
					STATUS_MIE <= 1'b0;
					STATUS_MPP <= PrivilegeModeW;
				end
				else if (P[1487]) begin
					STATUS_SPIE <= STATUS_SIE;
					STATUS_SIE <= 1'b0;
					STATUS_SPP <= PrivilegeModeW[0];
				end
			end
			else if (mretM) begin
				STATUS_MIE <= STATUS_MPIE;
				STATUS_MPIE <= 1'b1;
				STATUS_MPP <= (P[1486] ? P[1738-:2] : P[1742-:2]);
				STATUS_MPRV_INT <= STATUS_MPRV_INT & (STATUS_MPP == P[1742-:2]);
			end
			else if (sretM & P[1487]) begin
				STATUS_SIE <= STATUS_SPIE;
				STATUS_SPIE <= P[1487];
				STATUS_SPP <= 1'b0;
				STATUS_MPRV_INT <= 1'b0;
			end
			else if (WriteMSTATUSM) begin
				STATUS_TSR_INT <= P[1487] & CSRWriteValM[22];
				STATUS_TW_INT <= P[1486] & CSRWriteValM[21];
				STATUS_TVM_INT <= P[1487] & CSRWriteValM[20];
				STATUS_MXR_INT <= P[1487] & CSRWriteValM[19];
				STATUS_SUM_INT <= P[4067] & CSRWriteValM[18];
				STATUS_MPRV_INT <= P[1486] & CSRWriteValM[17];
				STATUS_FS_INT <= CSRWriteValM[14:13];
				STATUS_MPP <= STATUS_MPP_NEXT;
				STATUS_SPP <= P[1487] & CSRWriteValM[8];
				STATUS_MPIE <= CSRWriteValM[7];
				STATUS_SPIE <= P[1487] & CSRWriteValM[5];
				STATUS_MIE <= CSRWriteValM[3];
				STATUS_SIE <= P[1487] & CSRWriteValM[1];
				STATUS_UBE <= (P[1486] & P[4065]) & CSRWriteValM[6];
				STATUS_MBE <= nextMBE;
				STATUS_SBE <= nextSBE;
			end
			else if (($signed(P[4216-:32]) == 32) & WriteMSTATUSHM) begin
				STATUS_MBE <= P[4065] & CSRWriteValM[5];
				STATUS_SBE <= (P[1487] & P[4065]) & CSRWriteValM[4];
			end
			else if (P[1487] & WriteSSTATUSM) begin
				STATUS_MXR_INT <= P[1487] & CSRWriteValM[19];
				STATUS_SUM_INT <= P[4067] & CSRWriteValM[18];
				STATUS_FS_INT <= CSRWriteValM[14:13];
				STATUS_SPP <= P[1487] & CSRWriteValM[8];
				STATUS_SPIE <= P[1487] & CSRWriteValM[5];
				STATUS_SIE <= P[1487] & CSRWriteValM[1];
				STATUS_UBE <= (P[1486] & P[4065]) & CSRWriteValM[6];
			end
			else if ((FRegWriteM | WriteFRMM) | SetOrWriteFFLAGSM)
				STATUS_FS_INT <= 2'b11;
		end
	initial _sv2v_0 = 0;
endmodule
module csru (
	clk,
	reset,
	InstrValidNotFlushedM,
	CSRUWriteM,
	CSRAdrM,
	CSRWriteValM,
	STATUS_FS,
	CSRUReadValM,
	SetFflagsM,
	FRM_REGW,
	WriteFRMM,
	SetOrWriteFFLAGSM,
	IllegalCSRUAccessM
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire InstrValidNotFlushedM;
	input wire CSRUWriteM;
	input wire [11:0] CSRAdrM;
	input wire [$signed(P[4216-:32]) - 1:0] CSRWriteValM;
	input wire [1:0] STATUS_FS;
	output reg [$signed(P[4216-:32]) - 1:0] CSRUReadValM;
	input wire [4:0] SetFflagsM;
	output wire [2:0] FRM_REGW;
	output wire WriteFRMM;
	output wire SetOrWriteFFLAGSM;
	output reg IllegalCSRUAccessM;
	localparam FFLAGS = 12'h001;
	localparam FRM = 12'h002;
	localparam FCSR = 12'h003;
	wire [4:0] FFLAGS_REGW;
	wire [2:0] NextFRMM;
	wire [4:0] NextFFLAGSM;
	wire WriteFFLAGSM;
	assign WriteFRMM = (CSRUWriteM & (STATUS_FS != 2'b00)) & ((CSRAdrM == FRM) | (CSRAdrM == FCSR));
	assign WriteFFLAGSM = (CSRUWriteM & (STATUS_FS != 2'b00)) & ((CSRAdrM == FFLAGS) | (CSRAdrM == FCSR));
	assign NextFRMM = (CSRAdrM == FCSR ? CSRWriteValM[7:5] : CSRWriteValM[2:0]);
	assign NextFFLAGSM = (WriteFFLAGSM ? CSRWriteValM[4:0] : FFLAGS_REGW | SetFflagsM);
	assign SetOrWriteFFLAGSM = WriteFFLAGSM | (|SetFflagsM & InstrValidNotFlushedM);
	flopenr #(.WIDTH(3)) FRMreg(
		.clk(clk),
		.reset(reset),
		.en(WriteFRMM),
		.d(NextFRMM),
		.q(FRM_REGW)
	);
	flopenr #(.WIDTH(5)) FFLAGSreg(
		.clk(clk),
		.reset(reset),
		.en(SetOrWriteFFLAGSM),
		.d(NextFFLAGSM),
		.q(FFLAGS_REGW)
	);
	always @(*) begin
		if (_sv2v_0)
			;
		if (STATUS_FS == 2'b00) begin
			IllegalCSRUAccessM = 1'b1;
			CSRUReadValM = 1'sb0;
		end
		else begin
			IllegalCSRUAccessM = 1'b0;
			case (CSRAdrM)
				FFLAGS: CSRUReadValM = {{$signed(P[4216-:32]) - 5 {1'b0}}, FFLAGS_REGW};
				FRM: CSRUReadValM = {{$signed(P[4216-:32]) - 3 {1'b0}}, FRM_REGW};
				FCSR: CSRUReadValM = {{$signed(P[4216-:32]) - 8 {1'b0}}, FRM_REGW, FFLAGS_REGW};
				default: begin
					CSRUReadValM = 1'sb0;
					IllegalCSRUAccessM = 1'b1;
				end
			endcase
		end
	end
	initial _sv2v_0 = 0;
endmodule
module privdec (
	clk,
	reset,
	StallW,
	FlushW,
	InstrM,
	PrivilegedM,
	IllegalIEUFPUInstrM,
	IllegalCSRAccessM,
	PrivilegeModeW,
	STATUS_TSR,
	STATUS_TVM,
	STATUS_TW,
	IllegalInstrFaultM,
	EcallFaultM,
	BreakpointFaultM,
	sretM,
	mretM,
	RetM,
	wfiM,
	wfiW,
	sfencevmaM
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallW;
	input wire FlushW;
	input wire [31:15] InstrM;
	input wire PrivilegedM;
	input wire IllegalIEUFPUInstrM;
	input wire IllegalCSRAccessM;
	input wire [1:0] PrivilegeModeW;
	input wire STATUS_TSR;
	input wire STATUS_TVM;
	input wire STATUS_TW;
	output wire IllegalInstrFaultM;
	output wire EcallFaultM;
	output wire BreakpointFaultM;
	output wire sretM;
	output wire mretM;
	output wire RetM;
	output wire wfiM;
	output wire wfiW;
	output wire sfencevmaM;
	wire rs1zeroM;
	wire IllegalPrivilegedInstrM;
	wire WFITimeoutM;
	wire ebreakM;
	wire ecallM;
	wire sinvalvmaM;
	wire sfencewinvalM;
	wire sfenceinvalirM;
	wire invalM;
	assign rs1zeroM = InstrM[19:15] == 5'b00000;
	assign sinvalvmaM = InstrM[31:25] == 7'b0001011;
	assign sfencewinvalM = (InstrM[31:20] == 12'b000110000000) & rs1zeroM;
	assign sfenceinvalirM = (InstrM[31:20] == 12'b000110000001) & rs1zeroM;
	assign invalM = P[4055] & ((sinvalvmaM | sfencewinvalM) | sfenceinvalirM);
	assign sretM = (((PrivilegedM & (InstrM[31:20] == 12'b000100000010)) & rs1zeroM) & P[1487]) & ((PrivilegeModeW == P[1742-:2]) | ((PrivilegeModeW == P[1740-:2]) & ~STATUS_TSR));
	assign mretM = ((PrivilegedM & (InstrM[31:20] == 12'b001100000010)) & rs1zeroM) & (PrivilegeModeW == P[1742-:2]);
	assign RetM = sretM | mretM;
	assign ecallM = (PrivilegedM & (InstrM[31:20] == 12'b000000000000)) & rs1zeroM;
	assign ebreakM = (PrivilegedM & (InstrM[31:20] == 12'b000000000001)) & rs1zeroM;
	assign wfiM = (PrivilegedM & (InstrM[31:20] == 12'b000100000101)) & rs1zeroM;
	assign sfencevmaM = ((PrivilegedM & ((InstrM[31:25] == 7'b0001001) | invalM)) & ((PrivilegeModeW == P[1742-:2]) | ((PrivilegeModeW == P[1740-:2]) & ~STATUS_TVM))) & P[4067];
	generate
		if (P[1486]) begin : wfi
			wire [$signed(P[3632-:32]):0] WFICount;
			wire [$signed(P[3632-:32]):0] WFICountPlus1;
			assign WFICountPlus1 = (wfiM ? WFICount + 1 : {($signed(P[3632-:32]) >= 0 ? $signed(P[3632-:32]) + 1 : 1 - $signed(P[3632-:32])) {1'sb0}});
			flopr #(.WIDTH($signed(P[3632-:32]) + 1)) wficountreg(
				.clk(clk),
				.reset(reset),
				.d(WFICountPlus1),
				.q(WFICount)
			);
			assign WFITimeoutM = ((STATUS_TW & (PrivilegeModeW != P[1742-:2])) | (P[1487] & (PrivilegeModeW == P[1738-:2]))) & WFICount[$signed(P[3632-:32])];
		end
		else begin : genblk1
			assign WFITimeoutM = 1'b0;
		end
	endgenerate
	flopenrc #(.WIDTH(1)) wfiWReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(wfiM),
		.q(wfiW)
	);
	assign BreakpointFaultM = ebreakM;
	assign EcallFaultM = ecallM;
	assign IllegalPrivilegedInstrM = PrivilegedM & ~(((((sretM | mretM) | ecallM) | ebreakM) | wfiM) | sfencevmaM);
	assign IllegalInstrFaultM = ((IllegalIEUFPUInstrM | IllegalPrivilegedInstrM) | IllegalCSRAccessM) | WFITimeoutM;
endmodule
module privileged (
	clk,
	reset,
	StallD,
	StallE,
	StallM,
	StallW,
	FlushD,
	FlushE,
	FlushM,
	FlushW,
	CSRReadM,
	CSRWriteM,
	SrcAM,
	InstrM,
	InstrOrigM,
	IEUAdrxTvalM,
	PCM,
	InstrValidM,
	CommittedM,
	CommittedF,
	PrivilegedM,
	FRegWriteM,
	LoadStallD,
	StoreStallD,
	ICacheStallF,
	DCacheStallM,
	BPDirWrongM,
	BTAWrongM,
	RASPredPCWrongM,
	IClassWrongM,
	BPWrongM,
	IClassM,
	DCacheMiss,
	DCacheAccess,
	ICacheMiss,
	ICacheAccess,
	DivBusyE,
	FDivBusyE,
	InstrAccessFaultF,
	LoadAccessFaultM,
	StoreAmoAccessFaultM,
	HPTWInstrAccessFaultF,
	HPTWInstrPageFaultF,
	InstrPageFaultF,
	LoadPageFaultM,
	StoreAmoPageFaultM,
	InstrMisalignedFaultM,
	LoadMisalignedFaultM,
	StoreAmoMisalignedFaultM,
	IllegalIEUFPUInstrD,
	MTimerInt,
	MExtInt,
	SExtInt,
	MSwInt,
	MTIME_CLINT,
	SetFflagsM,
	SelHPTW,
	CSRReadValW,
	PrivilegeModeW,
	SATP_REGW,
	STATUS_MXR,
	STATUS_SUM,
	STATUS_MPRV,
	STATUS_MPP,
	STATUS_FS,
	PMPCFG_ARRAY_REGW,
	PMPADDR_ARRAY_REGW,
	FRM_REGW,
	ENVCFG_CBE,
	ENVCFG_PBMTE,
	ENVCFG_ADUE,
	EPCM,
	TrapVectorM,
	RetM,
	TrapM,
	sfencevmaM,
	InvalidateICacheM,
	BigEndianM,
	wfiM,
	IntPendingM
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallD;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushD;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	input wire CSRReadM;
	input wire CSRWriteM;
	input wire [$signed(P[4216-:32]) - 1:0] SrcAM;
	input wire [31:0] InstrM;
	input wire [31:0] InstrOrigM;
	input wire [$signed(P[4216-:32]) - 1:0] IEUAdrxTvalM;
	input wire [$signed(P[4216-:32]) - 1:0] PCM;
	input wire InstrValidM;
	input wire CommittedM;
	input wire CommittedF;
	input wire PrivilegedM;
	input wire FRegWriteM;
	input wire LoadStallD;
	input wire StoreStallD;
	input wire ICacheStallF;
	input wire DCacheStallM;
	input wire BPDirWrongM;
	input wire BTAWrongM;
	input wire RASPredPCWrongM;
	input wire IClassWrongM;
	input wire BPWrongM;
	input wire [3:0] IClassM;
	input wire DCacheMiss;
	input wire DCacheAccess;
	input wire ICacheMiss;
	input wire ICacheAccess;
	input wire DivBusyE;
	input wire FDivBusyE;
	input wire InstrAccessFaultF;
	input wire LoadAccessFaultM;
	input wire StoreAmoAccessFaultM;
	input wire HPTWInstrAccessFaultF;
	input wire HPTWInstrPageFaultF;
	input wire InstrPageFaultF;
	input wire LoadPageFaultM;
	input wire StoreAmoPageFaultM;
	input wire InstrMisalignedFaultM;
	input wire LoadMisalignedFaultM;
	input wire StoreAmoMisalignedFaultM;
	input wire IllegalIEUFPUInstrD;
	input wire MTimerInt;
	input wire MExtInt;
	input wire SExtInt;
	input wire MSwInt;
	input wire [63:0] MTIME_CLINT;
	input wire [4:0] SetFflagsM;
	input wire SelHPTW;
	output wire [$signed(P[4216-:32]) - 1:0] CSRReadValW;
	output wire [1:0] PrivilegeModeW;
	output wire [$signed(P[4216-:32]) - 1:0] SATP_REGW;
	output wire STATUS_MXR;
	output wire STATUS_SUM;
	output wire STATUS_MPRV;
	output wire [1:0] STATUS_MPP;
	output wire [1:0] STATUS_FS;
	output wire [($signed(P[3728-:32]) * 8) - 1:0] PMPCFG_ARRAY_REGW;
	output wire [(($signed(P[1640-:32]) - 3) >= 0 ? ($signed(P[3728-:32]) * ($signed(P[1640-:32]) - 2)) - 1 : ($signed(P[3728-:32]) * (4 - $signed(P[1640-:32]))) + ($signed(P[1640-:32]) - 4)):(($signed(P[1640-:32]) - 3) >= 0 ? 0 : $signed(P[1640-:32]) - 3)] PMPADDR_ARRAY_REGW;
	output wire [2:0] FRM_REGW;
	output wire [3:0] ENVCFG_CBE;
	output wire ENVCFG_PBMTE;
	output wire ENVCFG_ADUE;
	output wire [$signed(P[4216-:32]) - 1:0] EPCM;
	output wire [$signed(P[4216-:32]) - 1:0] TrapVectorM;
	output wire RetM;
	output wire TrapM;
	output wire sfencevmaM;
	input wire InvalidateICacheM;
	output wire BigEndianM;
	output wire wfiM;
	output wire IntPendingM;
	wire [3:0] CauseM;
	wire [15:0] MEDELEG_REGW;
	wire [11:0] MIDELEG_REGW;
	wire sretM;
	wire mretM;
	wire IllegalCSRAccessM;
	wire IllegalIEUFPUInstrM;
	wire InstrPageFaultM;
	wire InstrAccessFaultM;
	wire IllegalInstrFaultM;
	wire STATUS_SPP;
	wire STATUS_TSR;
	wire STATUS_TW;
	wire STATUS_TVM;
	wire STATUS_MIE;
	wire STATUS_SIE;
	wire [11:0] MIP_REGW;
	wire [11:0] MIE_REGW;
	wire [1:0] NextPrivilegeModeM;
	wire DelegateM;
	wire InterruptM;
	wire ExceptionM;
	wire HPTWInstrAccessFaultM;
	wire HPTWInstrPageFaultM;
	wire BreakpointFaultM;
	wire EcallFaultM;
	wire wfiW;
	privmode #(.P(P)) privmode(
		.clk(clk),
		.reset(reset),
		.StallW(StallW),
		.TrapM(TrapM),
		.mretM(mretM),
		.sretM(sretM),
		.DelegateM(DelegateM),
		.STATUS_MPP(STATUS_MPP),
		.STATUS_SPP(STATUS_SPP),
		.NextPrivilegeModeM(NextPrivilegeModeM),
		.PrivilegeModeW(PrivilegeModeW)
	);
	privdec #(.P(P)) pmd(
		.clk(clk),
		.reset(reset),
		.StallW(StallW),
		.FlushW(FlushW),
		.InstrM(InstrM[31:15]),
		.PrivilegedM(PrivilegedM),
		.IllegalIEUFPUInstrM(IllegalIEUFPUInstrM),
		.IllegalCSRAccessM(IllegalCSRAccessM),
		.PrivilegeModeW(PrivilegeModeW),
		.STATUS_TSR(STATUS_TSR),
		.STATUS_TVM(STATUS_TVM),
		.STATUS_TW(STATUS_TW),
		.IllegalInstrFaultM(IllegalInstrFaultM),
		.EcallFaultM(EcallFaultM),
		.BreakpointFaultM(BreakpointFaultM),
		.sretM(sretM),
		.mretM(mretM),
		.RetM(RetM),
		.wfiM(wfiM),
		.wfiW(wfiW),
		.sfencevmaM(sfencevmaM)
	);
	csr #(.P(P)) csr(
		.clk(clk),
		.reset(reset),
		.FlushM(FlushM),
		.FlushW(FlushW),
		.StallE(StallE),
		.StallM(StallM),
		.StallW(StallW),
		.InstrM(InstrM),
		.InstrOrigM(InstrOrigM),
		.PCM(PCM),
		.SrcAM(SrcAM),
		.IEUAdrxTvalM(IEUAdrxTvalM),
		.CSRReadM(CSRReadM),
		.CSRWriteM(CSRWriteM),
		.TrapM(TrapM),
		.mretM(mretM),
		.sretM(sretM),
		.InterruptM(InterruptM),
		.MTimerInt(MTimerInt),
		.MExtInt(MExtInt),
		.SExtInt(SExtInt),
		.MSwInt(MSwInt),
		.MTIME_CLINT(MTIME_CLINT),
		.InstrValidM(InstrValidM),
		.FRegWriteM(FRegWriteM),
		.LoadStallD(LoadStallD),
		.StoreStallD(StoreStallD),
		.BPDirWrongM(BPDirWrongM),
		.BTAWrongM(BTAWrongM),
		.RASPredPCWrongM(RASPredPCWrongM),
		.BPWrongM(BPWrongM),
		.sfencevmaM(sfencevmaM),
		.ExceptionM(ExceptionM),
		.InvalidateICacheM(InvalidateICacheM),
		.ICacheStallF(ICacheStallF),
		.DCacheStallM(DCacheStallM),
		.DivBusyE(DivBusyE),
		.FDivBusyE(FDivBusyE),
		.IClassWrongM(IClassWrongM),
		.IClassM(IClassM),
		.DCacheMiss(DCacheMiss),
		.DCacheAccess(DCacheAccess),
		.ICacheMiss(ICacheMiss),
		.ICacheAccess(ICacheAccess),
		.NextPrivilegeModeM(NextPrivilegeModeM),
		.PrivilegeModeW(PrivilegeModeW),
		.CauseM(CauseM),
		.SelHPTW(SelHPTW),
		.STATUS_MPP(STATUS_MPP),
		.STATUS_SPP(STATUS_SPP),
		.STATUS_TSR(STATUS_TSR),
		.STATUS_TVM(STATUS_TVM),
		.STATUS_MIE(STATUS_MIE),
		.STATUS_SIE(STATUS_SIE),
		.STATUS_MXR(STATUS_MXR),
		.STATUS_SUM(STATUS_SUM),
		.STATUS_MPRV(STATUS_MPRV),
		.STATUS_TW(STATUS_TW),
		.STATUS_FS(STATUS_FS),
		.MEDELEG_REGW(MEDELEG_REGW),
		.MIP_REGW(MIP_REGW),
		.MIE_REGW(MIE_REGW),
		.MIDELEG_REGW(MIDELEG_REGW),
		.SATP_REGW(SATP_REGW),
		.PMPCFG_ARRAY_REGW(PMPCFG_ARRAY_REGW),
		.PMPADDR_ARRAY_REGW(PMPADDR_ARRAY_REGW),
		.SetFflagsM(SetFflagsM),
		.FRM_REGW(FRM_REGW),
		.ENVCFG_CBE(ENVCFG_CBE),
		.ENVCFG_PBMTE(ENVCFG_PBMTE),
		.ENVCFG_ADUE(ENVCFG_ADUE),
		.EPCM(EPCM),
		.TrapVectorM(TrapVectorM),
		.CSRReadValW(CSRReadValW),
		.IllegalCSRAccessM(IllegalCSRAccessM),
		.BigEndianM(BigEndianM)
	);
	privpiperegs ppr(
		.clk(clk),
		.reset(reset),
		.StallD(StallD),
		.StallE(StallE),
		.StallM(StallM),
		.FlushD(FlushD),
		.FlushE(FlushE),
		.FlushM(FlushM),
		.InstrPageFaultF(InstrPageFaultF),
		.InstrAccessFaultF(InstrAccessFaultF),
		.HPTWInstrAccessFaultF(HPTWInstrAccessFaultF),
		.HPTWInstrPageFaultF(HPTWInstrPageFaultF),
		.IllegalIEUFPUInstrD(IllegalIEUFPUInstrD),
		.InstrPageFaultM(InstrPageFaultM),
		.InstrAccessFaultM(InstrAccessFaultM),
		.HPTWInstrAccessFaultM(HPTWInstrAccessFaultM),
		.HPTWInstrPageFaultM(HPTWInstrPageFaultM),
		.IllegalIEUFPUInstrM(IllegalIEUFPUInstrM)
	);
	trap #(.P(P)) trap(
		.reset(reset),
		.InstrMisalignedFaultM(InstrMisalignedFaultM),
		.InstrAccessFaultM(InstrAccessFaultM),
		.HPTWInstrAccessFaultM(HPTWInstrAccessFaultM),
		.HPTWInstrPageFaultM(HPTWInstrPageFaultM),
		.IllegalInstrFaultM(IllegalInstrFaultM),
		.BreakpointFaultM(BreakpointFaultM),
		.LoadMisalignedFaultM(LoadMisalignedFaultM),
		.StoreAmoMisalignedFaultM(StoreAmoMisalignedFaultM),
		.LoadAccessFaultM(LoadAccessFaultM),
		.StoreAmoAccessFaultM(StoreAmoAccessFaultM),
		.EcallFaultM(EcallFaultM),
		.InstrPageFaultM(InstrPageFaultM),
		.LoadPageFaultM(LoadPageFaultM),
		.StoreAmoPageFaultM(StoreAmoPageFaultM),
		.PrivilegeModeW(PrivilegeModeW),
		.MIP_REGW(MIP_REGW),
		.MIE_REGW(MIE_REGW),
		.MIDELEG_REGW(MIDELEG_REGW),
		.MEDELEG_REGW(MEDELEG_REGW),
		.STATUS_MIE(STATUS_MIE),
		.STATUS_SIE(STATUS_SIE),
		.InstrValidM(InstrValidM),
		.CommittedM(CommittedM),
		.CommittedF(CommittedF),
		.TrapM(TrapM),
		.wfiM(wfiM),
		.wfiW(wfiW),
		.InterruptM(InterruptM),
		.ExceptionM(ExceptionM),
		.IntPendingM(IntPendingM),
		.DelegateM(DelegateM),
		.CauseM(CauseM)
	);
endmodule
module privmode (
	clk,
	reset,
	StallW,
	TrapM,
	mretM,
	sretM,
	DelegateM,
	STATUS_MPP,
	STATUS_SPP,
	NextPrivilegeModeM,
	PrivilegeModeW
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallW;
	input wire TrapM;
	input wire mretM;
	input wire sretM;
	input wire DelegateM;
	input wire [1:0] STATUS_MPP;
	input wire STATUS_SPP;
	output reg [1:0] NextPrivilegeModeM;
	output wire [1:0] PrivilegeModeW;
	generate
		if (P[1486]) begin : privmode
			always @(*) begin
				if (_sv2v_0)
					;
				if (TrapM) begin
					if (P[1487] & DelegateM)
						NextPrivilegeModeM = P[1740-:2];
					else
						NextPrivilegeModeM = P[1742-:2];
				end
				else if (mretM)
					NextPrivilegeModeM = STATUS_MPP;
				else if (sretM)
					NextPrivilegeModeM = {1'b0, STATUS_SPP};
				else
					NextPrivilegeModeM = PrivilegeModeW;
			end
			flopenl #(.WIDTH(2)) privmodereg(
				.clk(clk),
				.load(reset),
				.en(~StallW),
				.d(NextPrivilegeModeM),
				.val(P[1742-:2]),
				.q(PrivilegeModeW)
			);
		end
		else begin : genblk1
			wire [2:1] sv2v_tmp_525FC;
			assign sv2v_tmp_525FC = P[1742-:2];
			always @(*) NextPrivilegeModeM = sv2v_tmp_525FC;
			assign PrivilegeModeW = P[1742-:2];
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module privpiperegs (
	clk,
	reset,
	StallD,
	StallE,
	StallM,
	FlushD,
	FlushE,
	FlushM,
	InstrPageFaultF,
	InstrAccessFaultF,
	HPTWInstrAccessFaultF,
	HPTWInstrPageFaultF,
	IllegalIEUFPUInstrD,
	InstrPageFaultM,
	InstrAccessFaultM,
	IllegalIEUFPUInstrM,
	HPTWInstrAccessFaultM,
	HPTWInstrPageFaultM
);
	input wire clk;
	input wire reset;
	input wire StallD;
	input wire StallE;
	input wire StallM;
	input wire FlushD;
	input wire FlushE;
	input wire FlushM;
	input wire InstrPageFaultF;
	input wire InstrAccessFaultF;
	input wire HPTWInstrAccessFaultF;
	input wire HPTWInstrPageFaultF;
	input wire IllegalIEUFPUInstrD;
	output wire InstrPageFaultM;
	output wire InstrAccessFaultM;
	output wire IllegalIEUFPUInstrM;
	output wire HPTWInstrAccessFaultM;
	output wire HPTWInstrPageFaultM;
	wire InstrPageFaultD;
	wire InstrAccessFaultD;
	wire HPTWInstrAccessFaultD;
	wire HPTWInstrPageFaultD;
	wire InstrPageFaultE;
	wire InstrAccessFaultE;
	wire HPTWInstrAccessFaultE;
	wire HPTWInstrPageFaultE;
	wire IllegalIEUFPUInstrE;
	flopenrc #(.WIDTH(4)) faultregD(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallD),
		.d({InstrPageFaultF, InstrAccessFaultF, HPTWInstrAccessFaultF, HPTWInstrPageFaultF}),
		.q({InstrPageFaultD, InstrAccessFaultD, HPTWInstrAccessFaultD, HPTWInstrPageFaultD})
	);
	flopenrc #(.WIDTH(5)) faultregE(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d({IllegalIEUFPUInstrD, InstrPageFaultD, InstrAccessFaultD, HPTWInstrAccessFaultD, HPTWInstrPageFaultD}),
		.q({IllegalIEUFPUInstrE, InstrPageFaultE, InstrAccessFaultE, HPTWInstrAccessFaultE, HPTWInstrPageFaultE})
	);
	flopenrc #(.WIDTH(5)) faultregM(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d({IllegalIEUFPUInstrE, InstrPageFaultE, InstrAccessFaultE, HPTWInstrAccessFaultE, HPTWInstrPageFaultE}),
		.q({IllegalIEUFPUInstrM, InstrPageFaultM, InstrAccessFaultM, HPTWInstrAccessFaultM, HPTWInstrPageFaultM})
	);
endmodule
module trap (
	reset,
	InstrMisalignedFaultM,
	InstrAccessFaultM,
	HPTWInstrAccessFaultM,
	HPTWInstrPageFaultM,
	IllegalInstrFaultM,
	BreakpointFaultM,
	LoadMisalignedFaultM,
	StoreAmoMisalignedFaultM,
	LoadAccessFaultM,
	StoreAmoAccessFaultM,
	EcallFaultM,
	InstrPageFaultM,
	LoadPageFaultM,
	StoreAmoPageFaultM,
	wfiM,
	wfiW,
	PrivilegeModeW,
	MIP_REGW,
	MIE_REGW,
	MIDELEG_REGW,
	MEDELEG_REGW,
	STATUS_MIE,
	STATUS_SIE,
	InstrValidM,
	CommittedM,
	CommittedF,
	TrapM,
	InterruptM,
	ExceptionM,
	IntPendingM,
	DelegateM,
	CauseM
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire reset;
	input wire InstrMisalignedFaultM;
	input wire InstrAccessFaultM;
	input wire HPTWInstrAccessFaultM;
	input wire HPTWInstrPageFaultM;
	input wire IllegalInstrFaultM;
	input wire BreakpointFaultM;
	input wire LoadMisalignedFaultM;
	input wire StoreAmoMisalignedFaultM;
	input wire LoadAccessFaultM;
	input wire StoreAmoAccessFaultM;
	input wire EcallFaultM;
	input wire InstrPageFaultM;
	input wire LoadPageFaultM;
	input wire StoreAmoPageFaultM;
	input wire wfiM;
	input wire wfiW;
	input wire [1:0] PrivilegeModeW;
	input wire [11:0] MIP_REGW;
	input wire [11:0] MIE_REGW;
	input wire [11:0] MIDELEG_REGW;
	input wire [15:0] MEDELEG_REGW;
	input wire STATUS_MIE;
	input wire STATUS_SIE;
	input wire InstrValidM;
	input wire CommittedM;
	input wire CommittedF;
	output wire TrapM;
	output wire InterruptM;
	output wire ExceptionM;
	output wire IntPendingM;
	output wire DelegateM;
	output reg [3:0] CauseM;
	wire MIntGlobalEnM;
	wire SIntGlobalEnM;
	wire Committed;
	wire BothInstrAccessFaultM;
	wire BothInstrPageFaultM;
	wire [11:0] PendingIntsM;
	wire [11:0] ValidIntsM;
	wire [11:0] EnabledIntsM;
	assign MIntGlobalEnM = (PrivilegeModeW != P[1742-:2]) | STATUS_MIE;
	assign SIntGlobalEnM = (PrivilegeModeW == P[1738-:2]) | ((PrivilegeModeW == P[1740-:2]) & STATUS_SIE);
	assign PendingIntsM = MIP_REGW & MIE_REGW;
	assign IntPendingM = |PendingIntsM;
	assign Committed = CommittedM | CommittedF;
	assign EnabledIntsM = (MIntGlobalEnM ? PendingIntsM & ~MIDELEG_REGW : {12 {1'sb0}}) | (SIntGlobalEnM ? PendingIntsM & MIDELEG_REGW : {12 {1'sb0}});
	assign ValidIntsM = (Committed ? {12 {1'sb0}} : EnabledIntsM);
	assign InterruptM = (|ValidIntsM & InstrValidM) & (~wfiM | wfiW);
	assign DelegateM = (P[1487] & (InterruptM ? MIDELEG_REGW[CauseM] : MEDELEG_REGW[CauseM])) & ((PrivilegeModeW == P[1738-:2]) | (PrivilegeModeW == P[1740-:2]));
	assign BothInstrAccessFaultM = InstrAccessFaultM | HPTWInstrAccessFaultM;
	assign BothInstrPageFaultM = InstrPageFaultM | HPTWInstrPageFaultM;
	assign ExceptionM = ((((((((((InstrMisalignedFaultM | BothInstrAccessFaultM) | IllegalInstrFaultM) | LoadMisalignedFaultM) | StoreAmoMisalignedFaultM) | BothInstrPageFaultM) | LoadPageFaultM) | StoreAmoPageFaultM) | BreakpointFaultM) | EcallFaultM) | LoadAccessFaultM) | StoreAmoAccessFaultM;
	assign TrapM = (ExceptionM & ~CommittedF) | InterruptM;
	always @(*) begin
		if (_sv2v_0)
			;
		if (reset)
			CauseM = 4'd0;
		else if (ValidIntsM[11])
			CauseM = 4'd11;
		else if (ValidIntsM[3])
			CauseM = 4'd3;
		else if (ValidIntsM[7])
			CauseM = 4'd7;
		else if (ValidIntsM[9])
			CauseM = 4'd9;
		else if (ValidIntsM[1])
			CauseM = 4'd1;
		else if (ValidIntsM[5])
			CauseM = 4'd5;
		else if (BothInstrPageFaultM)
			CauseM = 4'd12;
		else if (BothInstrAccessFaultM)
			CauseM = 4'd1;
		else if (IllegalInstrFaultM)
			CauseM = 4'd2;
		else if (InstrMisalignedFaultM)
			CauseM = 4'd0;
		else if (BreakpointFaultM)
			CauseM = 4'd3;
		else if (EcallFaultM)
			CauseM = {2'b10, PrivilegeModeW};
		else if (StoreAmoMisalignedFaultM & ~P[4059])
			CauseM = 4'd6;
		else if (LoadMisalignedFaultM & ~P[4059])
			CauseM = 4'd4;
		else if (StoreAmoPageFaultM)
			CauseM = 4'd15;
		else if (LoadPageFaultM)
			CauseM = 4'd13;
		else if (StoreAmoAccessFaultM)
			CauseM = 4'd7;
		else if (LoadAccessFaultM)
			CauseM = 4'd5;
		else if (StoreAmoMisalignedFaultM & P[4059])
			CauseM = 4'd6;
		else if (LoadMisalignedFaultM & P[4059])
			CauseM = 4'd4;
		else
			CauseM = 4'd0;
	end
	initial _sv2v_0 = 0;
endmodule
module csrindextoaddr (
	CSRWen,
	CSRAddr
);
	reg _sv2v_0;
	parameter TOTAL_CSRS = 36;
	input wire [TOTAL_CSRS - 1:0] CSRWen;
	output reg [11:0] CSRAddr;
	always @(*) begin
		if (_sv2v_0)
			;
		case (CSRWen)
			36'h000000000: CSRAddr = 12'h000;
			36'h000000001: CSRAddr = 12'h300;
			36'h000000002: CSRAddr = 12'h310;
			36'h000000004: CSRAddr = 12'h305;
			36'h000000008: CSRAddr = 12'h341;
			36'h000000010: CSRAddr = 12'h306;
			36'h000000020: CSRAddr = 12'h320;
			36'h000000040: CSRAddr = 12'h302;
			36'h000000080: CSRAddr = 12'h303;
			36'h000000100: CSRAddr = 12'h344;
			36'h000000200: CSRAddr = 12'h304;
			36'h000000400: CSRAddr = 12'h301;
			36'h000000800: CSRAddr = 12'h30a;
			36'h000001000: CSRAddr = 12'hf14;
			36'h000002000: CSRAddr = 12'h340;
			36'h000004000: CSRAddr = 12'h342;
			36'h000008000: CSRAddr = 12'h343;
			36'h000010000: CSRAddr = 12'hf11;
			36'h000020000: CSRAddr = 12'hf12;
			36'h000040000: CSRAddr = 12'hf13;
			36'h000080000: CSRAddr = 12'hf15;
			36'h000100000: CSRAddr = 12'h34a;
			36'h000200000: CSRAddr = 12'h100;
			36'h000400000: CSRAddr = 12'h104;
			36'h000800000: CSRAddr = 12'h105;
			36'h001000000: CSRAddr = 12'h141;
			36'h002000000: CSRAddr = 12'h106;
			36'h004000000: CSRAddr = 12'h10a;
			36'h008000000: CSRAddr = 12'h180;
			36'h010000000: CSRAddr = 12'h140;
			36'h020000000: CSRAddr = 12'h143;
			36'h040000000: CSRAddr = 12'h142;
			36'h080000000: CSRAddr = 12'h144;
			36'h100000000: CSRAddr = 12'h14d;
			36'h200000000: CSRAddr = 12'h001;
			36'h400000000: CSRAddr = 12'h002;
			36'h800000000: CSRAddr = 12'h003;
			default: CSRAddr = 12'h000;
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
module packetizer (
	rvvi,
	valid,
	m_axi_aclk,
	m_axi_aresetn,
	RVVIStall,
	RvviAxiWdata,
	RvviAxiWstrb,
	RvviAxiWlast,
	RvviAxiWvalid,
	RvviAxiWready
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter integer MAX_CSRS = 0;
	parameter [31:0] RVVI_INIT_TIME_OUT = 32'd4;
	parameter [31:0] RVVI_PACKET_DELAY = 32'd2;
	input wire [((72 + (5 * $signed(P[4216-:32]))) + (MAX_CSRS * ($signed(P[4216-:32]) + 16))) - 1:0] rvvi;
	input wire valid;
	input wire m_axi_aclk;
	input wire m_axi_aresetn;
	output wire RVVIStall;
	output wire [31:0] RvviAxiWdata;
	output wire [3:0] RvviAxiWstrb;
	output wire RvviAxiWlast;
	output wire RvviAxiWvalid;
	input wire RvviAxiWready;
	localparam NearTotalFrameLengthBits = (184 + (5 * $signed(P[4216-:32]))) + (MAX_CSRS * ($signed(P[4216-:32]) + 16));
	localparam WordPadLen = 32 - (NearTotalFrameLengthBits % 32);
	localparam TotalFrameLengthBits = NearTotalFrameLengthBits + WordPadLen;
	localparam TotalFrameLengthBytes = TotalFrameLengthBits / 8;
	wire [9:0] WordCount;
	wire [11:0] BytesInFrame;
	wire TransReady;
	wire BurstDone;
	wire WordCountReset;
	wire WordCountEnable;
	wire [47:0] SrcMac;
	wire [47:0] DstMac;
	wire [15:0] EthType;
	wire [15:0] Length;
	wire [TotalFrameLengthBits - 1:0] TotalFrame;
	wire [31:0] TotalFrameWords [(TotalFrameLengthBytes / 4) - 1:0];
	wire [WordPadLen - 1:0] WordPad;
	wire [((72 + (5 * $signed(P[4216-:32]))) + (MAX_CSRS * ($signed(P[4216-:32]) + 16))) - 1:0] rvviDelay;
	(* mark_debug = "true" *) reg [2:0] CurrState;
	(* mark_debug = "true" *) reg [2:0] NextState;
	wire [31:0] RstCount;
	(* mark_debug = "true" *) wire [31:0] FrameCount;
	wire RstCountRst;
	wire RstCountEn;
	wire CountFlag;
	wire DelayFlag;
	always @(posedge m_axi_aclk)
		if (~m_axi_aresetn)
			CurrState <= 3'd0;
		else
			CurrState <= NextState;
	always @(*) begin
		if (_sv2v_0)
			;
		case (CurrState)
			3'd0: NextState = 3'd1;
			3'd1:
				if (CountFlag)
					NextState = 3'd2;
				else
					NextState = 3'd1;
			3'd2:
				if (TransReady & valid)
					NextState = 3'd4;
				else if (~TransReady & valid)
					NextState = 3'd3;
				else
					NextState = 3'd2;
			3'd3:
				if (TransReady)
					NextState = 3'd4;
				else
					NextState = 3'd3;
			3'd4:
				if (BurstDone & TransReady)
					NextState = 3'd5;
				else
					NextState = 3'd4;
			3'd5:
				if (DelayFlag)
					NextState = 3'd2;
				else
					NextState = 3'd5;
			default: NextState = 3'd2;
		endcase
	end
	assign RVVIStall = CurrState != 3'd2;
	assign TransReady = RvviAxiWready;
	assign WordCountEnable = ((CurrState == 3'd2) & valid) | ((CurrState == 3'd4) & TransReady);
	assign WordCountReset = CurrState == 3'd2;
	assign RstCountEn = (CurrState == 3'd1) | (CurrState == 3'd5);
	assign RstCountRst = (CurrState == 3'd0) | (CurrState == 3'd4);
	counter #(.WIDTH(32)) rstcounter(
		.clk(m_axi_aclk),
		.reset(RstCountRst),
		.en(RstCountEn),
		.q(RstCount)
	);
	assign CountFlag = RstCount == RVVI_INIT_TIME_OUT;
	assign DelayFlag = RstCount == RVVI_PACKET_DELAY;
	counter #(.WIDTH(32)) framecounter(
		.clk(m_axi_aclk),
		.reset(~m_axi_aresetn),
		.en(RvviAxiWready & RvviAxiWlast),
		.q(FrameCount)
	);
	flopenr #(.WIDTH((72 + (5 * $signed(P[4216-:32]))) + (MAX_CSRS * ($signed(P[4216-:32]) + 16)))) rvvireg(
		.clk(m_axi_aclk),
		.reset(~m_axi_aresetn),
		.en(valid),
		.d(rvvi),
		.q(rvviDelay)
	);
	counter #(.WIDTH(10)) WordCounter(
		.clk(m_axi_aclk),
		.reset(WordCountReset),
		.en(WordCountEnable),
		.q(WordCount)
	);
	assign BytesInFrame = ((12'd2 + 12'd76) + (12'd6 + 12'd6)) + 12'd2;
	assign BurstDone = WordCount == (BytesInFrame[11:2] - 1'b1);
	genvar _gv_index_5;
	generate
		for (_gv_index_5 = 0; _gv_index_5 < (TotalFrameLengthBytes / 4); _gv_index_5 = _gv_index_5 + 1) begin : genblk1
			localparam index = _gv_index_5;
			assign TotalFrameWords[index] = TotalFrame[(index * 32) + 31:index * 32];
		end
	endgenerate
	assign Length = {4'b0000, BytesInFrame};
	assign WordPad = 1'sb0;
	assign TotalFrame = {WordPad, rvviDelay, EthType, DstMac, SrcMac};
	assign DstMac = 48'h8f5400001654;
	assign SrcMac = 48'h450211116843;
	assign EthType = 16'h005c;
	assign RvviAxiWdata = TotalFrameWords[WordCount[4:0]];
	assign RvviAxiWstrb = 1'sb1;
	assign RvviAxiWlast = BurstDone & (CurrState == 3'd4);
	assign RvviAxiWvalid = CurrState == 3'd4;
	initial _sv2v_0 = 0;
endmodule
module priorityaomux (
	Sel,
	A,
	Y,
	SelPriority
);
	parameter ROWS = 8;
	parameter COLS = 64;
	input wire [ROWS - 1:0] Sel;
	input wire [(ROWS * COLS) - 1:0] A;
	output wire [COLS - 1:0] Y;
	output wire [ROWS - 1:0] SelPriority;
	wire [(ROWS * COLS) - 1:0] AMasked;
	genvar _gv_index_6;
	priorityonehot #(.N(ROWS)) priorityonehot(
		.a(Sel),
		.y(SelPriority)
	);
	generate
		for (_gv_index_6 = 0; _gv_index_6 < ROWS; _gv_index_6 = _gv_index_6 + 1) begin : genblk1
			localparam index = _gv_index_6;
			assign AMasked[index * COLS+:COLS] = (SelPriority[index] ? A[index * COLS+:COLS] : {COLS * 1 {1'sb0}});
		end
	endgenerate
	or_rows #(
		.ROWS(ROWS),
		.COLS(COLS)
	) or_rows(
		.a(AMasked),
		.y(Y)
	);
endmodule
module regchangedetect (
	clk,
	reset,
	Value,
	Change
);
	parameter XLEN = 64;
	input clk;
	input reset;
	input wire [XLEN - 1:0] Value;
	output wire Change;
	wire [XLEN - 1:0] ValueD;
	flopr #(.WIDTH(XLEN)) register(
		.clk(clk),
		.reset(reset),
		.d(Value),
		.q(ValueD)
	);
	assign Change = |(Value ^ ValueD);
endmodule
module rvvisynth (
	clk,
	reset,
	StallE,
	StallM,
	StallW,
	FlushE,
	FlushM,
	FlushW,
	PCM,
	InstrValidM,
	InstrRawD,
	Mcycle,
	Minstret,
	TrapM,
	PrivilegeModeW,
	GPRWen,
	FPRWen,
	GPRAddr,
	FPRAddr,
	GPRValue,
	FPRValue,
	CSRArray,
	valid,
	rvvi
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter integer MAX_CSRS = 5;
	parameter integer TOTAL_CSRS = 36;
	input wire clk;
	input wire reset;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	input wire [$signed(P[4216-:32]) - 1:0] PCM;
	input wire InstrValidM;
	input wire [31:0] InstrRawD;
	input wire [63:0] Mcycle;
	input wire [63:0] Minstret;
	input wire TrapM;
	input wire [1:0] PrivilegeModeW;
	input wire GPRWen;
	input wire FPRWen;
	input wire [4:0] GPRAddr;
	input wire [4:0] FPRAddr;
	input wire [$signed(P[4216-:32]) - 1:0] GPRValue;
	input wire [$signed(P[4216-:32]) - 1:0] FPRValue;
	input wire [(TOTAL_CSRS * $signed(P[4216-:32])) - 1:0] CSRArray;
	output wire valid;
	output wire [((72 + (5 * $signed(P[4216-:32]))) + (MAX_CSRS * ($signed(P[4216-:32]) + 16))) - 1:0] rvvi;
	wire [$signed(P[4216-:32]) - 1:0] PCW;
	wire InstrValidW;
	wire [31:0] InstrRawE;
	wire [31:0] InstrRawM;
	wire [31:0] InstrRawW;
	wire TrapW;
	wire [$signed(P[4216-:32]) - 1:0] XLENZeros;
	wire [TOTAL_CSRS - 1:0] CSRArrayWen;
	wire [$signed(P[4216-:32]) - 1:0] CSRValue [MAX_CSRS - 1:0];
	wire [TOTAL_CSRS - 1:0] CSRWen [MAX_CSRS - 1:0];
	wire [11:0] CSRAddr [MAX_CSRS - 1:0];
	wire [MAX_CSRS - 1:0] EnabledCSRs;
	reg [MAX_CSRS - 1:0] CSRCountShort;
	wire [11:0] CSRCount;
	wire [(56 + (3 * $signed(P[4216-:32]))) - 1:0] Required;
	wire [(16 + (2 * $signed(P[4216-:32]))) - 1:0] Registers;
	wire [(MAX_CSRS * ($signed(P[4216-:32]) + 16)) - 1:0] CSRs;
	assign XLENZeros = 1'sb0;
	flopenrc #(.WIDTH(1)) InstrValidMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(InstrValidM),
		.q(InstrValidW)
	);
	flopenrc #(.WIDTH($signed(P[4216-:32]))) PCWReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(PCM),
		.q(PCW)
	);
	flopenrc #(.WIDTH(32)) InstrRawEReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(InstrRawD),
		.q(InstrRawE)
	);
	flopenrc #(.WIDTH(32)) InstrRawMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(InstrRawE),
		.q(InstrRawM)
	);
	flopenrc #(.WIDTH(32)) InstrRawWReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(InstrRawM),
		.q(InstrRawW)
	);
	flopenrc #(.WIDTH(1)) TrapWReg(
		.clk(clk),
		.reset(reset),
		.clear(1'b0),
		.en(~StallW),
		.d(TrapM),
		.q(TrapW)
	);
	assign valid = InstrValidW & ~StallW;
	assign Required = {4'b0000, CSRCount, 3'b000, FPRWen, GPRWen, PrivilegeModeW, TrapW, Minstret, Mcycle, InstrRawW, PCW};
	assign Registers = ({FPRWen, GPRWen} == 2'b11 ? {FPRValue, 3'b000, FPRAddr, GPRValue, 3'b000, GPRAddr} : ({FPRWen, GPRWen} == 2'b01 ? {XLENZeros, 8'b00000000, GPRValue, 3'b000, GPRAddr} : ({FPRWen, GPRWen} == 2'b10 ? {FPRValue, 3'b000, FPRAddr, XLENZeros, 8'b00000000} : {16 + (2 * $signed(P[4216-:32])) {1'sb0}})));
	genvar _gv_index_7;
	generate
		for (_gv_index_7 = 0; _gv_index_7 < TOTAL_CSRS; _gv_index_7 = _gv_index_7 + 1) begin : genblk1
			localparam index = _gv_index_7;
			regchangedetect #(.XLEN($signed(P[4216-:32]))) changedetect(
				.clk(clk),
				.reset(reset),
				.Value(CSRArray[index * $signed(P[4216-:32])+:$signed(P[4216-:32])]),
				.Change(CSRArrayWen[index])
			);
		end
	endgenerate
	wire [TOTAL_CSRS - 1:0] CSRWenPriorityMatrix [MAX_CSRS - 1:0];
	wire [TOTAL_CSRS - 1:0] CSRWenFilterMatrix [MAX_CSRS - 1:0];
	priorityaomux #(
		.ROWS(TOTAL_CSRS),
		.COLS($signed(P[4216-:32]))
	) firstpriorityaomux(
		.Sel(CSRArrayWen),
		.A(CSRArray),
		.Y(CSRValue[0]),
		.SelPriority(CSRWenPriorityMatrix[0])
	);
	assign CSRWenFilterMatrix[0] = CSRArrayWen;
	generate
		for (_gv_index_7 = 1; _gv_index_7 < MAX_CSRS; _gv_index_7 = _gv_index_7 + 1) begin : genblk2
			localparam index = _gv_index_7;
			priorityaomux #(
				.ROWS(TOTAL_CSRS),
				.COLS($signed(P[4216-:32]))
			) priorityaomux(
				.Sel(CSRWenFilterMatrix[index]),
				.A(CSRArray),
				.Y(CSRValue[index]),
				.SelPriority(CSRWenPriorityMatrix[index])
			);
			assign CSRWenFilterMatrix[index] = CSRWenFilterMatrix[index - 1] & ~CSRWenPriorityMatrix[index - 1];
		end
		for (_gv_index_7 = 0; _gv_index_7 < MAX_CSRS; _gv_index_7 = _gv_index_7 + 1) begin : genblk3
			localparam index = _gv_index_7;
			csrindextoaddr #(.TOTAL_CSRS(TOTAL_CSRS)) csrindextoaddr(
				.CSRWen(CSRWenPriorityMatrix[index]),
				.CSRAddr(CSRAddr[index])
			);
			assign CSRs[((index + 1) * ($signed(P[4216-:32]) + 16)) - 1:index * ($signed(P[4216-:32]) + 16)] = {CSRValue[index], 4'b0000, CSRAddr[index]};
			assign EnabledCSRs[index] = |CSRWenPriorityMatrix[index];
		end
	endgenerate
	integer index2;
	always @(*) begin
		if (_sv2v_0)
			;
		CSRCountShort = 1'sb0;
		for (index2 = 0; index2 < MAX_CSRS; index2 = index2 + 1)
			CSRCountShort = CSRCountShort + EnabledCSRs[index2];
	end
	assign CSRCount = {{{12 - MAX_CSRS} {1'b0}}, CSRCountShort};
	assign rvvi = {CSRs, Registers, Required};
	initial _sv2v_0 = 0;
endmodule
module triggergen (
	clk,
	reset,
	RvviAxiRdata,
	RvviAxiRstrb,
	RvviAxiRlast,
	RvviAxiRvalid,
	IlaTrigger
);
	reg _sv2v_0;
	input wire clk;
	input wire reset;
	input wire [31:0] RvviAxiRdata;
	input wire [3:0] RvviAxiRstrb;
	input wire RvviAxiRlast;
	input wire RvviAxiRvalid;
	output wire IlaTrigger;
	(* mark_debug = "true" *) reg [2:0] CurrState;
	(* mark_debug = "true" *) reg [2:0] NextState;
	wire [31:0] mem [4:0];
	wire [2:0] Counter;
	wire CounterEn;
	wire CounterRst;
	wire [31:0] RvviAxiRdataDelay;
	wire [3:0] RvviAxiRstrbDelay;
	wire RvviAxiRvalidDelay;
	wire Match;
	wire Overflow;
	wire Mismatch;
	wire Threshold;
	wire IlaTriggerOneCycle;
	assign mem[0] = 32'h11116843;
	assign mem[1] = 32'h16544502;
	assign mem[2] = 32'h8f540000;
	assign mem[3] = 32'h7274005c;
	assign mem[4] = 32'h6e696769;
	flopenr #(.WIDTH(32)) rvviaxirdatareg(
		.clk(clk),
		.reset(reset),
		.en(RvviAxiRvalid),
		.d(RvviAxiRdata),
		.q(RvviAxiRdataDelay)
	);
	flopenr #(.WIDTH(4)) rvviaxirstrbreg(
		.clk(clk),
		.reset(reset),
		.en(RvviAxiRvalid),
		.d(RvviAxiRstrb),
		.q(RvviAxiRstrbDelay)
	);
	flopr #(.WIDTH(1)) rvviaxirvalidreg(
		.clk(clk),
		.reset(reset),
		.d(RvviAxiRvalid),
		.q(RvviAxiRvalidDelay)
	);
	counter #(.WIDTH(3)) counter(
		.clk(clk),
		.reset(CounterRst),
		.en(CounterEn),
		.q(Counter)
	);
	always @(posedge clk)
		if (reset)
			CurrState <= 3'd0;
		else
			CurrState <= NextState;
	always @(*) begin
		if (_sv2v_0)
			;
		case (CurrState)
			3'd0:
				if (RvviAxiRvalid)
					NextState = 3'd1;
				else
					NextState = 3'd0;
			3'd1:
				if (RvviAxiRlast)
					NextState = 3'd0;
				else if (Mismatch | Overflow)
					NextState = 3'd2;
				else if (Threshold & Match)
					NextState = 3'd3;
				else
					NextState = 3'd1;
			3'd2:
				if (RvviAxiRlast)
					NextState = 3'd0;
				else
					NextState = 3'd2;
			3'd3:
				if (RvviAxiRlast)
					NextState = 3'd0;
				else
					NextState = 3'd4;
			3'd4:
				if (RvviAxiRlast)
					NextState = 3'd0;
				else
					NextState = 3'd4;
			default: NextState = 3'd0;
		endcase
	end
	assign Match = ((mem[Counter] == RvviAxiRdataDelay) & (CurrState == 3'd1)) & RvviAxiRvalidDelay;
	assign Overflow = Counter > 4'd4;
	assign Threshold = Counter >= 4'd4;
	assign Mismatch = ((mem[Counter] != RvviAxiRdataDelay) & (CurrState == 3'd1)) & RvviAxiRvalidDelay;
	assign IlaTriggerOneCycle = CurrState == 3'd3;
	assign CounterRst = CurrState == 3'd0;
	assign CounterEn = RvviAxiRvalid;
	wire [3:0] TriggerCount;
	wire TriggerReset;
	wire TriggerEn;
	counter #(.WIDTH(4)) triggercounter(
		.clk(clk),
		.reset(reset | TriggerReset),
		.en(TriggerEn),
		.q(TriggerCount)
	);
	assign TriggerReset = TriggerCount == 4'd10;
	assign TriggerEn = IlaTriggerOneCycle | ((TriggerCount != 4'd0) & (TriggerCount < 4'd10));
	assign IlaTrigger = TriggerEn;
	initial _sv2v_0 = 0;
endmodule
module ahbapbbridge (
	HCLK,
	HRESETn,
	HSEL,
	HADDR,
	HWDATA,
	HWSTRB,
	HWRITE,
	HTRANS,
	HREADY,
	HRDATA,
	HRESP,
	HREADYOUT,
	PCLK,
	PRESETn,
	PSEL,
	PWRITE,
	PENABLE,
	PADDR,
	PWDATA,
	PSTRB,
	PREADY,
	PRDATA
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter PERIPHS = 2;
	input wire HCLK;
	input wire HRESETn;
	input wire [PERIPHS - 1:0] HSEL;
	input wire [$signed(P[1640-:32]) - 1:0] HADDR;
	input wire [$signed(P[4216-:32]) - 1:0] HWDATA;
	input wire [($signed(P[4216-:32]) / 8) - 1:0] HWSTRB;
	input wire HWRITE;
	input wire [1:0] HTRANS;
	input wire HREADY;
	output reg [$signed(P[4216-:32]) - 1:0] HRDATA;
	output wire HRESP;
	output wire HREADYOUT;
	output wire PCLK;
	output wire PRESETn;
	output wire [PERIPHS - 1:0] PSEL;
	output wire PWRITE;
	output wire PENABLE;
	output wire [31:0] PADDR;
	output wire [$signed(P[4216-:32]) - 1:0] PWDATA;
	output wire [($signed(P[4216-:32]) / 8) - 1:0] PSTRB;
	input wire [PERIPHS - 1:0] PREADY;
	input wire [(PERIPHS * $signed(P[4216-:32])) - 1:0] PRDATA;
	wire initTrans;
	wire initTransSel;
	wire initTransSelD;
	wire nextPENABLE;
	reg PREADYOUT;
	assign PCLK = HCLK;
	assign PRESETn = HRESETn;
	assign initTrans = HTRANS[1] & HREADY;
	assign initTransSel = initTrans & |HSEL;
	flopen #(.WIDTH(32)) addrreg(
		.clk(HCLK),
		.en(HREADY),
		.d(HADDR[31:0]),
		.q(PADDR)
	);
	flopenr #(.WIDTH(1)) writereg(
		.clk(HCLK),
		.reset(~HRESETn),
		.en(HREADY),
		.d(HWRITE),
		.q(PWRITE)
	);
	flopenr #(.WIDTH(PERIPHS)) selreg(
		.clk(HCLK),
		.reset(~HRESETn),
		.en(HREADY),
		.d(HSEL & {PERIPHS {initTrans}}),
		.q(PSEL)
	);
	assign PWDATA = HWDATA;
	assign PSTRB = HWSTRB;
	flopr #(.WIDTH(1)) inittransreg(
		.clk(HCLK),
		.reset(~HRESETn),
		.d(initTransSel),
		.q(initTransSelD)
	);
	assign nextPENABLE = (PENABLE ? ~HREADY : initTransSelD);
	flopr #(.WIDTH(1)) enablereg(
		.clk(HCLK),
		.reset(~HRESETn),
		.d(nextPENABLE),
		.q(PENABLE)
	);
	reg signed [31:0] i;
	always @(*) begin
		if (_sv2v_0)
			;
		HRDATA = 1'sb0;
		PREADYOUT = 1'b1;
		for (i = 0; i < PERIPHS; i = i + 1)
			if (PSEL[i]) begin
				HRDATA = PRDATA[i * $signed(P[4216-:32])+:$signed(P[4216-:32])];
				PREADYOUT = PREADY[i];
			end
	end
	assign HREADYOUT = PREADYOUT & ~initTransSelD;
	assign HRESP = 1'b0;
	initial _sv2v_0 = 0;
endmodule
module clint_apb (
	PCLK,
	PRESETn,
	PSEL,
	PADDR,
	PWDATA,
	PSTRB,
	PWRITE,
	PENABLE,
	PRDATA,
	PREADY,
	MTIME,
	MTimerInt,
	MSwInt
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire PCLK;
	input wire PRESETn;
	input wire PSEL;
	input wire [15:0] PADDR;
	input wire [$signed(P[4216-:32]) - 1:0] PWDATA;
	input wire [($signed(P[4216-:32]) / 8) - 1:0] PSTRB;
	input wire PWRITE;
	input wire PENABLE;
	output reg [$signed(P[4216-:32]) - 1:0] PRDATA;
	output wire PREADY;
	output reg [63:0] MTIME;
	output wire MTimerInt;
	output wire MSwInt;
	localparam CLINT_MSIP = 16'h0000;
	localparam CLINT_MTIMECMP = 16'h4000;
	localparam CLINT_MTIME = 16'hbff8;
	reg MSIP;
	wire [15:0] entry;
	wire memwrite;
	reg [63:0] MTIMECMP;
	integer i;
	integer j;
	assign memwrite = (PWRITE & PENABLE) & PSEL;
	assign PREADY = 1'b1;
	generate
		if ($signed(P[4216-:32]) == 64) begin : genblk1
			assign entry = {PADDR[15:3], 3'b000};
		end
		else begin : genblk1
			assign entry = {PADDR[15:2], 2'b00};
		end
		if ($signed(P[4216-:32]) == 64) begin : clint
			always @(posedge PCLK)
				case (entry)
					CLINT_MSIP: PRDATA <= {63'b000000000000000000000000000000000000000000000000000000000000000, MSIP};
					CLINT_MTIMECMP: PRDATA <= MTIMECMP;
					CLINT_MTIME: PRDATA <= MTIME;
					default: PRDATA <= 1'sb0;
				endcase
			always @(posedge PCLK)
				if (~PRESETn) begin
					MSIP <= 1'b0;
					MTIMECMP <= 64'hffffffffffffffff;
				end
				else if (memwrite) begin
					if (entry == CLINT_MSIP)
						MSIP <= PWDATA[0];
					if (entry == CLINT_MTIMECMP) begin
						for (i = 0; i < ($signed(P[4216-:32]) / 8); i = i + 1)
							if (PSTRB[i])
								MTIMECMP[i * 8+:8] <= PWDATA[i * 8+:8];
					end
				end
			always @(posedge PCLK)
				if (~PRESETn)
					MTIME <= 1'sb0;
				else if (memwrite & (entry == 16'hbff8)) begin
					for (j = 0; j < ($signed(P[4216-:32]) / 8); j = j + 1)
						if (PSTRB[j])
							MTIME[j * 8+:8] <= PWDATA[j * 8+:8];
				end
				else
					MTIME <= MTIME + 1;
		end
		else begin : clint
			always @(posedge PCLK)
				case (entry)
					16'h0000: PRDATA <= {31'b0000000000000000000000000000000, MSIP};
					16'h4000: PRDATA <= MTIMECMP[31:0];
					16'h4004: PRDATA <= MTIMECMP[63:32];
					16'hbff8: PRDATA <= MTIME[31:0];
					16'hbffc: PRDATA <= MTIME[63:32];
					default: PRDATA <= 1'sb0;
				endcase
			always @(posedge PCLK)
				if (~PRESETn) begin
					MSIP <= 1'b0;
					MTIMECMP <= 64'hffffffffffffffff;
				end
				else if (memwrite) begin
					if (entry == 16'h0000)
						MSIP <= PWDATA[0];
					if (entry == 16'h4000) begin
						for (j = 0; j < ($signed(P[4216-:32]) / 8); j = j + 1)
							if (PSTRB[j])
								MTIMECMP[j * 8+:8] <= PWDATA[j * 8+:8];
					end
					if (entry == 16'h4004) begin
						for (j = 0; j < ($signed(P[4216-:32]) / 8); j = j + 1)
							if (PSTRB[j])
								MTIMECMP[32 + (j * 8)+:8] <= PWDATA[j * 8+:8];
					end
				end
			always @(posedge PCLK)
				if (~PRESETn)
					MTIME <= 1'sb0;
				else if (memwrite & (entry == 16'hbff8)) begin
					for (i = 0; i < ($signed(P[4216-:32]) / 8); i = i + 1)
						if (PSTRB[i])
							MTIME[i * 8+:8] <= PWDATA[i * 8+:8];
				end
				else if (memwrite & (entry == 16'hbffc)) begin
					for (i = 0; i < ($signed(P[4216-:32]) / 8); i = i + 1)
						if (PSTRB[i])
							MTIME[32 + (i * 8)+:8] <= PWDATA[i * 8+:8];
				end
				else
					MTIME <= MTIME + 1;
		end
	endgenerate
	assign MSwInt = MSIP;
	assign MTimerInt = {1'b0, MTIME} >= {1'b0, MTIMECMP};
endmodule
module gpio_apb (
	PCLK,
	PRESETn,
	PSEL,
	PADDR,
	PWDATA,
	PSTRB,
	PWRITE,
	PENABLE,
	PRDATA,
	PREADY,
	iof0,
	iof1,
	GPIOIN,
	GPIOOUT,
	GPIOEN,
	GPIOIntr
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire PCLK;
	input wire PRESETn;
	input wire PSEL;
	input wire [7:0] PADDR;
	input wire [$signed(P[4216-:32]) - 1:0] PWDATA;
	input wire [($signed(P[4216-:32]) / 8) - 1:0] PSTRB;
	input wire PWRITE;
	input wire PENABLE;
	output wire [$signed(P[4216-:32]) - 1:0] PRDATA;
	output wire PREADY;
	input wire [31:0] iof0;
	input wire [31:0] iof1;
	input wire [31:0] GPIOIN;
	output wire [31:0] GPIOOUT;
	output wire [31:0] GPIOEN;
	output wire GPIOIntr;
	localparam GPIO_INPUT_VAL = 8'h00;
	localparam GPIO_INPUT_EN = 8'h04;
	localparam GPIO_OUTPUT_EN = 8'h08;
	localparam GPIO_OUTPUT_VAL = 8'h0c;
	localparam GPIO_RISE_IE = 8'h18;
	localparam GPIO_RISE_IP = 8'h1c;
	localparam GPIO_FALL_IE = 8'h20;
	localparam GPIO_FALL_IP = 8'h24;
	localparam GPIO_HIGH_IE = 8'h28;
	localparam GPIO_HIGH_IP = 8'h2c;
	localparam GPIO_LOW_IE = 8'h30;
	localparam GPIO_LOW_IP = 8'h34;
	localparam GPIO_IOF_EN = 8'h38;
	localparam GPIO_IOF_SEL = 8'h3c;
	localparam GPIO_OUT_XOR = 8'h40;
	wire [31:0] input0d;
	wire [31:0] input1d;
	wire [31:0] input2d;
	wire [31:0] input3d;
	wire [31:0] input_val;
	reg [31:0] input_en;
	reg [31:0] output_en;
	reg [31:0] output_val;
	reg [31:0] rise_ie;
	reg [31:0] rise_ip;
	reg [31:0] fall_ie;
	reg [31:0] fall_ip;
	reg [31:0] high_ie;
	reg [31:0] high_ip;
	reg [31:0] low_ie;
	reg [31:0] low_ip;
	reg [31:0] out_xor;
	reg [31:0] iof_en;
	reg [31:0] iof_sel;
	wire [31:0] iof_out;
	wire [31:0] gpio_out;
	wire [7:0] entry;
	wire [31:0] Din;
	reg [31:0] Dout;
	wire memwrite;
	assign entry = {PADDR[7:2], 2'b00};
	assign memwrite = (PWRITE & PENABLE) & PSEL;
	assign PREADY = 1'b1;
	assign Din = PWDATA[31:0];
	generate
		if ($signed(P[4216-:32]) == 64) begin : genblk1
			assign PRDATA = {Dout, Dout};
		end
		else begin : genblk1
			assign PRDATA = Dout;
		end
	endgenerate
	always @(posedge PCLK)
		if (~PRESETn) begin
			input_en <= 1'sb0;
			output_en <= 1'sb0;
			output_val <= 1'sb0;
			rise_ie <= 1'sb0;
			rise_ip <= 1'sb0;
			fall_ie <= 1'sb0;
			fall_ip <= 1'sb0;
			high_ie <= 1'sb0;
			high_ip <= 1'sb0;
			low_ie <= 1'sb0;
			low_ip <= 1'sb0;
			iof_en <= 1'sb0;
			iof_sel <= 1'sb0;
			out_xor <= 1'sb0;
		end
		else begin
			if (memwrite)
				case (entry)
					GPIO_INPUT_EN: input_en <= Din;
					GPIO_OUTPUT_EN: output_en <= Din;
					GPIO_OUTPUT_VAL: output_val <= Din;
					GPIO_RISE_IE: rise_ie <= Din;
					GPIO_FALL_IE: fall_ie <= Din;
					GPIO_HIGH_IE: high_ie <= Din;
					GPIO_LOW_IE: low_ie <= Din;
					GPIO_IOF_EN: iof_en <= Din;
					GPIO_IOF_SEL: iof_sel <= Din;
					GPIO_OUT_XOR: out_xor <= Din;
				endcase
			if (memwrite & (entry == GPIO_RISE_IP))
				rise_ip <= rise_ip & ~Din;
			else
				rise_ip <= rise_ip | (input2d & ~input3d);
			if (memwrite & (entry == GPIO_FALL_IP))
				fall_ip <= fall_ip & ~Din;
			else
				fall_ip <= fall_ip | (~input2d & input3d);
			if (memwrite & (entry == GPIO_HIGH_IP))
				high_ip <= high_ip & ~Din;
			else
				high_ip <= high_ip | input3d;
			if (memwrite & (entry == GPIO_LOW_IP))
				low_ip <= low_ip & ~Din;
			else
				low_ip <= low_ip | ~input3d;
			case (entry)
				GPIO_INPUT_VAL: Dout <= input_val;
				GPIO_INPUT_EN: Dout <= input_en;
				GPIO_OUTPUT_EN: Dout <= output_en;
				GPIO_OUTPUT_VAL: Dout <= output_val;
				GPIO_RISE_IE: Dout <= rise_ie;
				GPIO_RISE_IP: Dout <= rise_ip;
				GPIO_FALL_IE: Dout <= fall_ie;
				GPIO_FALL_IP: Dout <= fall_ip;
				GPIO_HIGH_IE: Dout <= high_ie;
				GPIO_HIGH_IP: Dout <= high_ip;
				GPIO_LOW_IE: Dout <= low_ie;
				GPIO_LOW_IP: Dout <= low_ip;
				GPIO_IOF_EN: Dout <= iof_en;
				GPIO_IOF_SEL: Dout <= iof_sel;
				GPIO_OUT_XOR: Dout <= out_xor;
				default: Dout <= 1'sb0;
			endcase
		end
	generate
		if (P[2179]) begin : genblk2
			assign input0d = ((output_en & GPIOOUT) | (~output_en & GPIOIN)) & input_en;
		end
		else begin : genblk2
			assign input0d = GPIOIN & input_en;
		end
	endgenerate
	flop #(.WIDTH(32)) sync1(
		.clk(PCLK),
		.d(input0d),
		.q(input1d)
	);
	flop #(.WIDTH(32)) sync2(
		.clk(PCLK),
		.d(input1d),
		.q(input2d)
	);
	flop #(.WIDTH(32)) sync3(
		.clk(PCLK),
		.d(input2d),
		.q(input3d)
	);
	assign input_val = input3d;
	assign iof_out = (iof_sel & iof1) | (~iof_sel & iof0);
	assign gpio_out = (iof_en & iof_out) | (~iof_en & output_val);
	assign GPIOOUT = gpio_out ^ out_xor;
	assign GPIOEN = output_en;
	assign GPIOIntr = |{rise_ip & rise_ie, fall_ip & fall_ie, high_ip & high_ie, low_ip & low_ie};
endmodule
module plic_apb (
	PCLK,
	PRESETn,
	PSEL,
	PADDR,
	PWDATA,
	PSTRB,
	PWRITE,
	PENABLE,
	PRDATA,
	PREADY,
	UARTIntr,
	GPIOIntr,
	SPIIntr,
	SDCIntr,
	MExtInt,
	SExtInt
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire PCLK;
	input wire PRESETn;
	input wire PSEL;
	input wire [27:0] PADDR;
	input wire [$signed(P[4216-:32]) - 1:0] PWDATA;
	input wire [($signed(P[4216-:32]) / 8) - 1:0] PSTRB;
	input wire PWRITE;
	input wire PENABLE;
	output wire [$signed(P[4216-:32]) - 1:0] PRDATA;
	output wire PREADY;
	input wire UARTIntr;
	input wire GPIOIntr;
	input wire SPIIntr;
	input wire SDCIntr;
	output wire MExtInt;
	output wire SExtInt;
	localparam PLIC_INTPRIORITY0 = 24'h000000;
	localparam PLIC_INTPENDING0 = 24'h001000;
	localparam PLIC_INTPENDING1 = 24'h001004;
	localparam PLIC_INTEN00 = 24'h002000;
	localparam PLIC_INTEN01 = 24'h002004;
	localparam PLIC_INTEN10 = 24'h002080;
	localparam PLIC_INTEN11 = 24'h002084;
	localparam PLIC_THRESHOLD0 = 24'h200000;
	localparam PLIC_CLAIMCOMPLETE0 = 24'h200004;
	localparam PLIC_THRESHOLD1 = 24'h201000;
	localparam PLIC_CLAIMCOMPLETE1 = 24'h201004;
	wire memwrite;
	wire memread;
	wire [23:0] entry;
	wire [31:0] Din;
	reg [31:0] Dout;
	reg [$signed(P[2145-:32]):1] requests;
	reg [($signed(P[2145-:32]) >= 1 ? ($signed(P[2145-:32]) * 3) + 2 : ((2 - $signed(P[2145-:32])) * 3) + (($signed(P[2145-:32]) * 3) - 1)):($signed(P[2145-:32]) >= 1 ? 3 : $signed(P[2145-:32]) * 3)] intPriority;
	reg [$signed(P[2145-:32]):1] intInProgress;
	wire [$signed(P[2145-:32]):1] intPending;
	wire [$signed(P[2145-:32]):1] nextIntPending;
	reg [5:0] intThreshold;
	reg [($signed(P[2145-:32]) >= 1 ? (2 * $signed(P[2145-:32])) + 0 : (2 * (2 - $signed(P[2145-:32]))) + ($signed(P[2145-:32]) - 1)):($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32]) + 0)] intEn;
	reg [11:0] intClaim;
	wire [($signed(P[2145-:32]) >= 1 ? (14 * $signed(P[2145-:32])) + ((1 + $signed(P[2145-:32])) - 1) : (14 * (2 - $signed(P[2145-:32]))) + (($signed(P[2145-:32]) + (2 - $signed(P[2145-:32]))) - 1)):($signed(P[2145-:32]) >= 1 ? 1 + $signed(P[2145-:32]) : $signed(P[2145-:32]) + (2 - $signed(P[2145-:32])))] irqMatrix;
	wire [14:1] priorities_with_irqs;
	wire [14:1] max_priority_with_irqs;
	wire [($signed(P[2145-:32]) >= 1 ? (2 * $signed(P[2145-:32])) + 0 : (2 * (2 - $signed(P[2145-:32]))) + ($signed(P[2145-:32]) - 1)):($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32]) + 0)] irqs_at_max_priority;
	reg [14:1] threshMask;
	wire [$signed(P[2145-:32]) - 1:0] One;
	localparam PLIC_SRC_TOP = ($signed(P[2145-:32]) >= 32 ? $signed(P[2145-:32]) : 1);
	localparam PLIC_SRC_BOT = ($signed(P[2145-:32]) >= 32 ? 32 : 1);
	localparam PLIC_SRC_DINTOP = ($signed(P[2145-:32]) >= 32 ? $signed(P[2145-:32]) - 32 : 0);
	localparam PLIC_SRC_EXT = ($signed(P[2145-:32]) >= 32 ? 63 - $signed(P[2145-:32]) : 31);
	assign memwrite = (PWRITE & PENABLE) & PSEL;
	assign memread = ~PWRITE & PSEL;
	assign PREADY = 1'b1;
	assign entry = {PADDR[23:2], 2'b00};
	assign One[$signed(P[2145-:32]) - 1:1] = 1'sb0;
	assign One[0] = 1'b1;
	assign Din = PWDATA[31:0];
	generate
		if ($signed(P[4216-:32]) == 64) begin : genblk1
			assign PRDATA = {Dout, Dout};
		end
		else begin : genblk1
			assign PRDATA = Dout;
		end
	endgenerate
	localparam PLIC_NUM_SRC_MIN_32 = ($signed(P[2145-:32]) < 32 ? $signed(P[2145-:32]) : 31);
	always @(posedge PCLK)
		if (~PRESETn) begin
			intPriority <= 1'sb0;
			intEn <= 1'sb0;
			intThreshold <= 1'sb0;
			intInProgress <= 1'sb0;
		end
		else begin
			if (memwrite)
				casez (entry)
					24'h0000zz: intPriority[($signed(P[2145-:32]) >= 1 ? entry[7:2] : 1 - (entry[7:2] - $signed(P[2145-:32]))) * 3+:3] <= Din[2:0];
					PLIC_INTEN00: intEn[($signed(P[2145-:32]) >= 1 ? 0 + ($signed(P[2145-:32]) >= 1 ? (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) : 1 - ((PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) - $signed(P[2145-:32]))) : ((0 + ($signed(P[2145-:32]) >= 1 ? (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) : 1 - ((PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) - $signed(P[2145-:32])))) + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1)-:(PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)] <= Din[PLIC_NUM_SRC_MIN_32:1];
					PLIC_INTEN10: intEn[($signed(P[2145-:32]) >= 1 ? ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])) + ($signed(P[2145-:32]) >= 1 ? (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) : 1 - ((PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) - $signed(P[2145-:32]))) : ((($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])) + ($signed(P[2145-:32]) >= 1 ? (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) : 1 - ((PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) - $signed(P[2145-:32])))) + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1)-:(PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)] <= Din[PLIC_NUM_SRC_MIN_32:1];
					PLIC_INTEN01:
						if ($signed(P[2145-:32]) >= 32)
							intEn[($signed(P[2145-:32]) >= 1 ? 0 + ($signed(P[2145-:32]) >= 1 ? (PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) : 1 - ((PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) - $signed(P[2145-:32]))) : ((0 + ($signed(P[2145-:32]) >= 1 ? (PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) : 1 - ((PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) - $signed(P[2145-:32])))) + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1)-:(PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)] <= Din[PLIC_SRC_DINTOP:0];
					PLIC_INTEN11:
						if ($signed(P[2145-:32]) >= 32)
							intEn[($signed(P[2145-:32]) >= 1 ? ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])) + ($signed(P[2145-:32]) >= 1 ? (PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) : 1 - ((PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) - $signed(P[2145-:32]))) : ((($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])) + ($signed(P[2145-:32]) >= 1 ? (PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) : 1 - ((PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) - $signed(P[2145-:32])))) + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1)-:(PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)] <= Din[PLIC_SRC_DINTOP:0];
					PLIC_THRESHOLD0: intThreshold[0+:3] <= Din[2:0];
					PLIC_CLAIMCOMPLETE0: intInProgress <= intInProgress & ~(One << (Din[5:0] - 1));
					PLIC_THRESHOLD1: intThreshold[3+:3] <= Din[2:0];
					PLIC_CLAIMCOMPLETE1: intInProgress <= intInProgress & ~(One << (Din[5:0] - 1));
				endcase
			if (memread)
				casez (entry)
					PLIC_INTPRIORITY0: Dout <= 32'b00000000000000000000000000000000;
					24'h0000zz: Dout <= {29'b00000000000000000000000000000, intPriority[($signed(P[2145-:32]) >= 1 ? entry[7:2] : 1 - (entry[7:2] - $signed(P[2145-:32]))) * 3+:3]};
					PLIC_INTPENDING0: Dout <= {{31 - PLIC_NUM_SRC_MIN_32 {1'b0}}, intPending[PLIC_NUM_SRC_MIN_32:1], 1'b0};
					PLIC_INTEN00: Dout <= {{31 - PLIC_NUM_SRC_MIN_32 {1'b0}}, intEn[($signed(P[2145-:32]) >= 1 ? 0 + ($signed(P[2145-:32]) >= 1 ? (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) : 1 - ((PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) - $signed(P[2145-:32]))) : ((0 + ($signed(P[2145-:32]) >= 1 ? (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) : 1 - ((PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) - $signed(P[2145-:32])))) + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1)-:(PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)], 1'b0};
					PLIC_INTPENDING1:
						if ($signed(P[2145-:32]) >= 32)
							Dout <= {{PLIC_SRC_EXT {1'b0}}, intPending[PLIC_SRC_TOP:PLIC_SRC_BOT]};
					PLIC_INTEN01:
						if ($signed(P[2145-:32]) >= 32)
							Dout <= {{PLIC_SRC_EXT {1'b0}}, intEn[($signed(P[2145-:32]) >= 1 ? 0 + ($signed(P[2145-:32]) >= 1 ? (PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) : 1 - ((PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) - $signed(P[2145-:32]))) : ((0 + ($signed(P[2145-:32]) >= 1 ? (PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) : 1 - ((PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) - $signed(P[2145-:32])))) + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1)-:(PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)]};
					PLIC_INTEN10: Dout <= {{31 - PLIC_NUM_SRC_MIN_32 {1'b0}}, intEn[($signed(P[2145-:32]) >= 1 ? ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])) + ($signed(P[2145-:32]) >= 1 ? (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) : 1 - ((PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) - $signed(P[2145-:32]))) : ((($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])) + ($signed(P[2145-:32]) >= 1 ? (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) : 1 - ((PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : (PLIC_NUM_SRC_MIN_32 + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1) - $signed(P[2145-:32])))) + (PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)) - 1)-:(PLIC_NUM_SRC_MIN_32 >= 1 ? PLIC_NUM_SRC_MIN_32 : 2 - PLIC_NUM_SRC_MIN_32)], 1'b0};
					PLIC_INTEN11:
						if ($signed(P[2145-:32]) >= 32)
							Dout <= {{PLIC_SRC_EXT {1'b0}}, intEn[($signed(P[2145-:32]) >= 1 ? ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])) + ($signed(P[2145-:32]) >= 1 ? (PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) : 1 - ((PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) - $signed(P[2145-:32]))) : ((($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])) + ($signed(P[2145-:32]) >= 1 ? (PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) : 1 - ((PLIC_SRC_TOP >= PLIC_SRC_BOT ? PLIC_SRC_TOP : (PLIC_SRC_TOP + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1) - $signed(P[2145-:32])))) + (PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)) - 1)-:(PLIC_SRC_TOP >= PLIC_SRC_BOT ? (PLIC_SRC_TOP - PLIC_SRC_BOT) + 1 : (PLIC_SRC_BOT - PLIC_SRC_TOP) + 1)]};
					PLIC_THRESHOLD0: Dout <= {29'b00000000000000000000000000000, intThreshold[0+:3]};
					PLIC_CLAIMCOMPLETE0: begin
						Dout <= {26'b00000000000000000000000000, intClaim[0+:6]};
						intInProgress <= intInProgress | (One << (intClaim[0+:6] - 1));
					end
					PLIC_THRESHOLD1: Dout <= {29'b00000000000000000000000000000, intThreshold[3+:3]};
					PLIC_CLAIMCOMPLETE1: begin
						Dout <= {26'b00000000000000000000000000, intClaim[6+:6]};
						intInProgress <= intInProgress | (One << (intClaim[6+:6] - 1));
					end
					default: Dout <= 32'h00000000;
				endcase
			else
				Dout <= 32'h00000000;
		end
	always @(*) begin
		if (_sv2v_0)
			;
		requests = {$signed(P[2145-:32]) {1'b0}};
		if ($signed(P[2112-:32]) != 0)
			requests[$signed(P[2112-:32])] = GPIOIntr;
		if ($signed(P[2080-:32]) != 0)
			requests[$signed(P[2080-:32])] = UARTIntr;
		if ($signed(P[2048-:32]) != 0)
			requests[$signed(P[2048-:32])] = SPIIntr;
		if ($signed(P[2016-:32]) != 0)
			requests[$signed(P[2016-:32])] = SDCIntr;
	end
	assign nextIntPending = (intPending | requests) & ~intInProgress;
	flopr #(.WIDTH($signed(P[2145-:32]))) intPendingFlop(
		.clk(PCLK),
		.reset(~PRESETn),
		.d(nextIntPending),
		.q(intPending)
	);
	genvar _gv_ctx_1;
	generate
		for (_gv_ctx_1 = 0; _gv_ctx_1 < 2; _gv_ctx_1 = _gv_ctx_1 + 1) begin : genblk2
			localparam ctx = _gv_ctx_1;
			genvar _gv_src_1;
			genvar _gv_pri_1;
			for (_gv_pri_1 = 1; _gv_pri_1 <= 7; _gv_pri_1 = _gv_pri_1 + 1) begin : genblk1
				localparam pri = _gv_pri_1;
				for (_gv_src_1 = 1; _gv_src_1 <= $signed(P[2145-:32]); _gv_src_1 = _gv_src_1 + 1) begin : genblk1
					localparam src = _gv_src_1;
					assign irqMatrix[(((ctx * 7) + pri) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))) + ($signed(P[2145-:32]) >= 1 ? src : 1 - (src - $signed(P[2145-:32])))] = ((intPriority[($signed(P[2145-:32]) >= 1 ? src : 1 - (src - $signed(P[2145-:32]))) * 3+:3] == pri) & intPending[src]) & intEn[(ctx * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))) + ($signed(P[2145-:32]) >= 1 ? src : 1 - (src - $signed(P[2145-:32])))];
				end
			end
			assign priorities_with_irqs[(ctx * 7) + 7-:7] = {|irqMatrix[($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32])) + (((ctx * 7) + 7) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])))+:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))], |irqMatrix[($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32])) + (((ctx * 7) + 6) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])))+:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))], |irqMatrix[($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32])) + (((ctx * 7) + 5) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])))+:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))], |irqMatrix[($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32])) + (((ctx * 7) + 4) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])))+:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))], |irqMatrix[($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32])) + (((ctx * 7) + 3) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])))+:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))], |irqMatrix[($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32])) + (((ctx * 7) + 2) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])))+:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))], |irqMatrix[($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32])) + (((ctx * 7) + 1) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])))+:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))]};
			assign max_priority_with_irqs[(ctx * 7) + 7-:7] = {priorities_with_irqs[(ctx * 7) + 7], priorities_with_irqs[(ctx * 7) + 6] & ~|priorities_with_irqs[(ctx * 7) + 7], priorities_with_irqs[(ctx * 7) + 5] & ~|priorities_with_irqs[(ctx * 7) + 7-:2], priorities_with_irqs[(ctx * 7) + 4] & ~|priorities_with_irqs[(ctx * 7) + 7-:3], priorities_with_irqs[(ctx * 7) + 3] & ~|priorities_with_irqs[(ctx * 7) + 7-:4], priorities_with_irqs[(ctx * 7) + 2] & ~|priorities_with_irqs[(ctx * 7) + 7-:5], priorities_with_irqs[(ctx * 7) + 1] & ~|priorities_with_irqs[(ctx * 7) + 7-:6]};
			assign irqs_at_max_priority[($signed(P[2145-:32]) >= 1 ? (ctx * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))) + ($signed(P[2145-:32]) >= 1 ? ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : ($signed(P[2145-:32]) + ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))) - 1) : 1 - (($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : ($signed(P[2145-:32]) + ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))) - 1) - $signed(P[2145-:32]))) : (((ctx * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))) + ($signed(P[2145-:32]) >= 1 ? ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : ($signed(P[2145-:32]) + ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))) - 1) : 1 - (($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : ($signed(P[2145-:32]) + ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))) - 1) - $signed(P[2145-:32])))) + ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))) - 1)-:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))] = (((((({$signed(P[2145-:32]) {max_priority_with_irqs[(ctx * 7) + 7]}} & irqMatrix[($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32])) + (((ctx * 7) + 7) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])))+:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))]) | ({$signed(P[2145-:32]) {max_priority_with_irqs[(ctx * 7) + 6]}} & irqMatrix[($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32])) + (((ctx * 7) + 6) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])))+:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))])) | ({$signed(P[2145-:32]) {max_priority_with_irqs[(ctx * 7) + 5]}} & irqMatrix[($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32])) + (((ctx * 7) + 5) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])))+:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))])) | ({$signed(P[2145-:32]) {max_priority_with_irqs[(ctx * 7) + 4]}} & irqMatrix[($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32])) + (((ctx * 7) + 4) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])))+:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))])) | ({$signed(P[2145-:32]) {max_priority_with_irqs[(ctx * 7) + 3]}} & irqMatrix[($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32])) + (((ctx * 7) + 3) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])))+:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))])) | ({$signed(P[2145-:32]) {max_priority_with_irqs[(ctx * 7) + 2]}} & irqMatrix[($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32])) + (((ctx * 7) + 2) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])))+:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))])) | ({$signed(P[2145-:32]) {max_priority_with_irqs[(ctx * 7) + 1]}} & irqMatrix[($signed(P[2145-:32]) >= 1 ? 1 : $signed(P[2145-:32])) + (((ctx * 7) + 1) * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32])))+:($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))]);
			integer k;
			always @(*) begin
				if (_sv2v_0)
					;
				intClaim[ctx * 6+:6] = 6'b000000;
				for (k = $signed(P[2145-:32]); k > 0; k = k - 1)
					if (irqs_at_max_priority[(ctx * ($signed(P[2145-:32]) >= 1 ? $signed(P[2145-:32]) : 2 - $signed(P[2145-:32]))) + ($signed(P[2145-:32]) >= 1 ? k : 1 - (k - $signed(P[2145-:32])))])
						intClaim[ctx * 6+:6] = k[5:0];
			end
			always @(*) begin
				if (_sv2v_0)
					;
				threshMask[(ctx * 7) + 7] = intThreshold[ctx * 3+:3] != 7;
				threshMask[(ctx * 7) + 6] = (intThreshold[ctx * 3+:3] != 6) & threshMask[(ctx * 7) + 7];
				threshMask[(ctx * 7) + 5] = (intThreshold[ctx * 3+:3] != 5) & threshMask[(ctx * 7) + 6];
				threshMask[(ctx * 7) + 4] = (intThreshold[ctx * 3+:3] != 4) & threshMask[(ctx * 7) + 5];
				threshMask[(ctx * 7) + 3] = (intThreshold[ctx * 3+:3] != 3) & threshMask[(ctx * 7) + 4];
				threshMask[(ctx * 7) + 2] = (intThreshold[ctx * 3+:3] != 2) & threshMask[(ctx * 7) + 3];
				threshMask[(ctx * 7) + 1] = (intThreshold[ctx * 3+:3] != 1) & threshMask[(ctx * 7) + 2];
			end
		end
	endgenerate
	assign MExtInt = |(threshMask[1+:7] & priorities_with_irqs[1+:7]);
	assign SExtInt = |(threshMask[8+:7] & priorities_with_irqs[8+:7]);
	initial _sv2v_0 = 0;
endmodule
module ram_ahb (
	HCLK,
	HRESETn,
	HSELRam,
	HADDR,
	HWRITE,
	HREADY,
	HTRANS,
	HWDATA,
	HWSTRB,
	HREADRam,
	HRESPRam,
	HREADYRam
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter RANGE = 65535;
	parameter PRELOAD = 0;
	input wire HCLK;
	input wire HRESETn;
	input wire HSELRam;
	input wire [$signed(P[1640-:32]) - 1:0] HADDR;
	input wire HWRITE;
	input wire HREADY;
	input wire [1:0] HTRANS;
	input wire [$signed(P[4216-:32]) - 1:0] HWDATA;
	input wire [($signed(P[4216-:32]) / 8) - 1:0] HWSTRB;
	output wire [$signed(P[4216-:32]) - 1:0] HREADRam;
	output wire HRESPRam;
	output wire HREADYRam;
	localparam ADDR_WIDTH = $clog2(RANGE / 8);
	localparam OFFSET = $clog2($signed(P[4216-:32]) / 8);
	wire [($signed(P[4216-:32]) / 8) - 1:0] ByteMask;
	wire [$signed(P[1640-:32]) - 1:0] HADDRD;
	wire [$signed(P[1640-:32]) - 1:0] RamAddr;
	wire initTrans;
	wire memwrite;
	wire memwriteD;
	wire memread;
	wire nextHREADYRam;
	wire DelayReady;
	assign initTrans = (HREADY & HSELRam) & HTRANS[1];
	assign memwrite = initTrans & HWRITE;
	assign memread = initTrans & ~HWRITE;
	flopenr #(.WIDTH(1)) memwritereg(
		.clk(HCLK),
		.reset(~HRESETn),
		.en(HREADY),
		.d(memwrite),
		.q(memwriteD)
	);
	flopenr #(.WIDTH($signed(P[1640-:32]))) haddrreg(
		.clk(HCLK),
		.reset(~HRESETn),
		.en(HREADY),
		.d(HADDR),
		.q(HADDRD)
	);
	assign nextHREADYRam = ~(memwriteD & memread) & ~DelayReady;
	flopr #(.WIDTH(1)) readyreg(
		.clk(HCLK),
		.reset(~HRESETn),
		.d(nextHREADYRam),
		.q(HREADYRam)
	);
	assign HRESPRam = 1'b0;
	mux2 #(.WIDTH($signed(P[1640-:32]))) adrmux(
		.d0(HADDR),
		.d1(HADDRD),
		.s(memwriteD | ~HREADY),
		.y(RamAddr)
	);
	ram1p1rwbe #(
		.USE_SRAM(P[1743]),
		.DEPTH(RANGE / 8),
		.WIDTH($signed(P[4216-:32])),
		.PRELOAD_ENABLED(PRELOAD)
	) memory(
		.clk(HCLK),
		.ce(1'b1),
		.addr(RamAddr[(ADDR_WIDTH + OFFSET) - 1:OFFSET]),
		.we(memwriteD),
		.din(HWDATA),
		.bwe(HWSTRB),
		.dout(HREADRam)
	);
	generate
		if ($signed(P[4119-:32]) > 0) begin : genblk1
			wire [7:0] NextCycle;
			wire [7:0] Cycle;
			wire CntEn;
			wire CntRst;
			wire CycleFlag;
			flopenr #(.WIDTH(8)) counter(
				.clk(HCLK),
				.reset(~HRESETn | CntRst),
				.en(CntEn),
				.d(NextCycle),
				.q(Cycle)
			);
			assign NextCycle = Cycle + 1'b1;
			reg CurrState;
			reg NextState;
			always @(posedge HCLK)
				if (~HRESETn)
					CurrState <= 1'd0;
				else
					CurrState <= NextState;
			always @(*) begin
				if (_sv2v_0)
					;
				case (CurrState)
					1'd0:
						if (initTrans & ~CycleFlag)
							NextState = 1'd1;
						else
							NextState = 1'd0;
					1'd1:
						if (CycleFlag)
							NextState = 1'd0;
						else
							NextState = 1'd1;
					default: NextState = 1'd0;
				endcase
			end
			assign CycleFlag = Cycle == P[4095:4088];
			assign CntEn = NextState == 1'd1;
			assign DelayReady = NextState == 1'd1;
			assign CntRst = NextState == 1'd0;
		end
		else begin : genblk1
			assign DelayReady = 1'b0;
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module rom_ahb (
	HCLK,
	HRESETn,
	HSELRom,
	HADDR,
	HREADY,
	HTRANS,
	HREADRom,
	HRESPRom,
	HREADYRom
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter RANGE = 65535;
	parameter PRELOAD = 0;
	input wire HCLK;
	input wire HRESETn;
	input wire HSELRom;
	input wire [$signed(P[1640-:32]) - 1:0] HADDR;
	input wire HREADY;
	input wire [1:0] HTRANS;
	output wire [$signed(P[4216-:32]) - 1:0] HREADRom;
	output wire HRESPRom;
	output wire HREADYRom;
	localparam ADDR_WIDTH = $clog2(RANGE / 8);
	localparam OFFSET = $clog2($signed(P[4216-:32]) / 8);
	assign HREADYRom = 1'b1;
	assign HRESPRom = 1'b0;
	rom1p1r #(
		.ADDR_WIDTH(ADDR_WIDTH),
		.DATA_WIDTH($signed(P[4216-:32])),
		.PRELOAD_ENABLED(PRELOAD)
	) memory(
		.clk(HCLK),
		.ce(1'b1),
		.addr(HADDR[(ADDR_WIDTH + OFFSET) - 1:OFFSET]),
		.dout(HREADRom)
	);
endmodule
module spi_apb (
	PCLK,
	PRESETn,
	PSEL,
	PADDR,
	PWDATA,
	PSTRB,
	PWRITE,
	PENABLE,
	PREADY,
	PRDATA,
	SPIOut,
	SPIIn,
	SPICS,
	SPIIntr,
	SPICLK
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire PCLK;
	input wire PRESETn;
	input wire PSEL;
	input wire [7:0] PADDR;
	input wire [$signed(P[4216-:32]) - 1:0] PWDATA;
	input wire [($signed(P[4216-:32]) / 8) - 1:0] PSTRB;
	input wire PWRITE;
	input wire PENABLE;
	output wire PREADY;
	output wire [$signed(P[4216-:32]) - 1:0] PRDATA;
	output wire SPIOut;
	input wire SPIIn;
	output wire [3:0] SPICS;
	output wire SPIIntr;
	output wire SPICLK;
	localparam SPI_SCKDIV = 8'h00;
	localparam SPI_SCKMODE = 8'h04;
	localparam SPI_CSID = 8'h10;
	localparam SPI_CSDEF = 8'h14;
	localparam SPI_CSMODE = 8'h18;
	localparam SPI_DELAY0 = 8'h28;
	localparam SPI_DELAY1 = 8'h2c;
	localparam SPI_FMT = 8'h40;
	localparam SPI_TXDATA = 8'h48;
	localparam SPI_RXDATA = 8'h4c;
	localparam SPI_TXMARK = 8'h50;
	localparam SPI_RXMARK = 8'h54;
	localparam SPI_IE = 8'h70;
	localparam SPI_IP = 8'h74;
	reg [11:0] SckDiv;
	reg [1:0] SckMode;
	reg [1:0] ChipSelectID;
	reg [3:0] ChipSelectDef;
	reg [1:0] ChipSelectMode;
	reg [15:0] Delay0;
	reg [15:0] Delay1;
	reg [4:0] Format;
	wire [7:0] ReceiveData;
	reg [8:0] TransmitData;
	reg [2:0] TransmitWatermark;
	reg [2:0] ReceiveWatermark;
	reg [1:0] InterruptEnable;
	reg [1:0] InterruptPending;
	wire [7:0] Entry;
	wire Memwrite;
	wire [31:0] Din;
	reg [31:0] Dout;
	wire SCLKenable;
	wire EndOfFrame;
	wire Transmitting;
	wire InactiveState;
	wire [3:0] FrameLength;
	wire ResetSCLKenable;
	wire TransmitStart;
	reg TransmitStartD;
	reg [1:0] CurrState;
	reg [1:0] NextState;
	wire TransmitWriteMark;
	wire TransmitReadMark;
	wire ReceiveWriteMark;
	wire ReceiveReadMark;
	wire TransmitFIFOFull;
	wire TransmitFIFOEmpty;
	wire TransmitFIFOWriteInc;
	wire TransmitFIFOReadInc;
	wire [7:0] TransmitReadData;
	wire ReceiveFIFOWriteInc;
	wire ReceiveFIFOReadInc;
	wire ReceiveFIFOFull;
	wire ReceiveFIFOEmpty;
	wire [2:0] TransmitWriteWatermarkLevel;
	wire [2:0] ReceiveReadWatermarkLevel;
	wire [7:0] ReceiveShiftRegEndian;
	wire ShiftEdge;
	wire SampleEdge;
	reg [7:0] TransmitReg;
	reg [7:0] ReceiveShiftReg;
	wire [7:0] TransmitDataEndian;
	wire TransmitLoad;
	reg TransmitRegLoaded;
	wire ShiftIn;
	wire [3:0] LeftShiftAmount;
	wire [7:0] ASR;
	reg [3:0] ChipSelectAuto;
	wire [3:0] ChipSelectInternal;
	assign Entry = {PADDR[7:2], 2'b00};
	assign Memwrite = (PWRITE & PENABLE) & PSEL;
	assign PREADY = 1'b1;
	assign Din = PWDATA[31:0];
	generate
		if ($signed(P[4216-:32]) == 64) begin : genblk1
			assign PRDATA = {Dout, Dout};
		end
		else begin : genblk1
			assign PRDATA = Dout;
		end
	endgenerate
	always @(posedge PCLK)
		if (~PRESETn) begin
			SckDiv <= 12'd3;
			SckMode <= 2'b00;
			ChipSelectID <= 2'b00;
			ChipSelectDef <= 4'b1111;
			ChipSelectMode <= 2'b00;
			Delay0 <= 16'b0000000100000001;
			Delay1 <= 16'b0000000000000001;
			Format <= 5'b10000;
			TransmitData <= 9'b000000000;
			TransmitWatermark <= 3'b000;
			ReceiveWatermark <= 3'b000;
			InterruptEnable <= 2'b00;
			InterruptPending <= 2'b00;
		end
		else begin
			if (Memwrite)
				case (Entry)
					SPI_SCKDIV: SckDiv <= Din[11:0];
					SPI_SCKMODE: SckMode <= Din[1:0];
					SPI_CSID: ChipSelectID <= Din[1:0];
					SPI_CSDEF: ChipSelectDef <= Din[3:0];
					SPI_CSMODE: ChipSelectMode <= Din[1:0];
					SPI_DELAY0: Delay0 <= {Din[23:16], Din[7:0]};
					SPI_DELAY1: Delay1 <= {Din[23:16], Din[7:0]};
					SPI_FMT: Format <= {Din[19:16], Din[2]};
					SPI_TXDATA:
						if (~TransmitFIFOFull)
							TransmitData[7:0] <= Din[7:0];
					SPI_TXMARK: TransmitWatermark <= Din[2:0];
					SPI_RXMARK: ReceiveWatermark <= Din[2:0];
					SPI_IE: InterruptEnable <= Din[1:0];
				endcase
			InterruptPending[0] <= TransmitReadMark;
			InterruptPending[1] <= ReceiveWriteMark;
			case (Entry)
				SPI_SCKDIV: Dout <= {20'b00000000000000000000, SckDiv};
				SPI_SCKMODE: Dout <= {30'b000000000000000000000000000000, SckMode};
				SPI_CSID: Dout <= {30'b000000000000000000000000000000, ChipSelectID};
				SPI_CSDEF: Dout <= {28'b0000000000000000000000000000, ChipSelectDef};
				SPI_CSMODE: Dout <= {30'b000000000000000000000000000000, ChipSelectMode};
				SPI_DELAY0: Dout <= {8'b00000000, Delay0[15:8], 8'b00000000, Delay0[7:0]};
				SPI_DELAY1: Dout <= {8'b00000000, Delay1[15:8], 8'b00000000, Delay1[7:0]};
				SPI_FMT: Dout <= {12'b000000000000, Format[4:1], 13'b0000000000000, Format[0], 2'b00};
				SPI_TXDATA: Dout <= {TransmitFIFOFull, 31'b0000000000000000000000000000000};
				SPI_RXDATA: Dout <= {ReceiveFIFOEmpty, 23'b00000000000000000000000, ReceiveData[7:0]};
				SPI_TXMARK: Dout <= {29'b00000000000000000000000000000, TransmitWatermark};
				SPI_RXMARK: Dout <= {29'b00000000000000000000000000000, ReceiveWatermark};
				SPI_IE: Dout <= {30'b000000000000000000000000000000, InterruptEnable};
				SPI_IP: Dout <= {30'b000000000000000000000000000000, InterruptPending};
				default: Dout <= 32'b00000000000000000000000000000000;
			endcase
		end
	assign ResetSCLKenable = Memwrite & (Entry == SPI_SCKDIV);
	assign FrameLength = Format[4:1];
	spi_controller controller(
		.PCLK(PCLK),
		.PRESETn(PRESETn),
		.TransmitStart(TransmitStart),
		.TransmitRegLoaded(TransmitRegLoaded),
		.ResetSCLKenable(ResetSCLKenable),
		.SckDiv(SckDiv),
		.SckMode(SckMode),
		.CSMode(ChipSelectMode),
		.Delay0(Delay0),
		.Delay1(Delay1),
		.FrameLength(FrameLength),
		.TransmitFIFOEmpty(TransmitFIFOEmpty),
		.SCLKenable(SCLKenable),
		.ShiftEdge(ShiftEdge),
		.SampleEdge(SampleEdge),
		.EndOfFrame(EndOfFrame),
		.Transmitting(Transmitting),
		.InactiveState(InactiveState),
		.SPICLK(SPICLK)
	);
	flopr #(.WIDTH(1)) txwincreg(
		.clk(PCLK),
		.reset(~PRESETn),
		.d((Memwrite & (Entry == SPI_TXDATA)) & ~TransmitFIFOFull),
		.q(TransmitFIFOWriteInc)
	);
	flopenr #(.WIDTH(1)) txrincreg(
		.clk(PCLK),
		.reset(~PRESETn),
		.en(SCLKenable),
		.d(TransmitStartD | (EndOfFrame & ~TransmitFIFOEmpty)),
		.q(TransmitFIFOReadInc)
	);
	always @(posedge PCLK)
		if (~PRESETn)
			TransmitRegLoaded <= 1'b0;
		else if (TransmitLoad)
			TransmitRegLoaded <= 1'b1;
		else if (ShiftEdge | EndOfFrame)
			TransmitRegLoaded <= 1'b0;
	always @(posedge PCLK)
		if (~PRESETn)
			CurrState <= 2'd0;
		else
			CurrState <= NextState;
	always @(*) begin
		if (_sv2v_0)
			;
		case (CurrState)
			2'd0:
				if (~TransmitFIFOEmpty & ~Transmitting)
					NextState = 2'd1;
				else
					NextState = 2'd0;
			2'd1: NextState = 2'd2;
			2'd2:
				if (~Transmitting & ~TransmitRegLoaded)
					NextState = 2'd0;
				else
					NextState = 2'd2;
			default: NextState = 2'd0;
		endcase
	end
	assign TransmitStart = CurrState == 2'd1;
	always @(posedge PCLK)
		if (~PRESETn)
			TransmitStartD <= 1'b0;
		else if (TransmitStart)
			TransmitStartD <= 1'b1;
		else if (SCLKenable)
			TransmitStartD <= 1'b0;
	spi_fifo #(
		.M(3),
		.N(8)
	) txFIFO(
		.PCLK(PCLK),
		.wen(1'b1),
		.ren(SCLKenable),
		.PRESETn(PRESETn),
		.winc(TransmitFIFOWriteInc),
		.rinc(TransmitFIFOReadInc),
		.wdata(TransmitData[7:0]),
		.wwatermarklevel(TransmitWriteWatermarkLevel),
		.rwatermarklevel(TransmitWatermark[2:0]),
		.rdata(TransmitReadData[7:0]),
		.wfull(TransmitFIFOFull),
		.rempty(TransmitFIFOEmpty),
		.wwatermark(TransmitWriteMark),
		.rwatermark(TransmitReadMark)
	);
	flopr #(.WIDTH(1)) rxfiforincreg(
		.clk(PCLK),
		.reset(~PRESETn),
		.d((((Entry == SPI_RXDATA) & ~ReceiveFIFOEmpty) & PSEL) & ~ReceiveFIFOReadInc),
		.q(ReceiveFIFOReadInc)
	);
	flopenr #(.WIDTH(1)) rxfifowincreg(
		.clk(PCLK),
		.reset(~PRESETn),
		.en(SCLKenable),
		.d(EndOfFrame),
		.q(ReceiveFIFOWriteInc)
	);
	spi_fifo #(
		.M(3),
		.N(8)
	) rxFIFO(
		.PCLK(PCLK),
		.wen(SCLKenable),
		.ren(1'b1),
		.PRESETn(PRESETn),
		.winc(ReceiveFIFOWriteInc),
		.rinc(ReceiveFIFOReadInc),
		.wdata(ReceiveShiftRegEndian),
		.wwatermarklevel(ReceiveWatermark[2:0]),
		.rwatermarklevel(ReceiveReadWatermarkLevel),
		.rdata(ReceiveData[7:0]),
		.wfull(ReceiveFIFOFull),
		.rempty(ReceiveFIFOEmpty),
		.wwatermark(ReceiveWriteMark),
		.rwatermark(ReceiveReadMark)
	);
	assign TransmitLoad = TransmitStart | (EndOfFrame & ~TransmitFIFOEmpty);
	function automatic [7:0] _sv2v_strm_D90CD;
		input reg [7:0] inp;
		reg [7:0] _sv2v_strm_BEEC1_inp;
		reg [7:0] _sv2v_strm_BEEC1_out;
		integer _sv2v_strm_BEEC1_idx;
		begin
			_sv2v_strm_BEEC1_inp = {inp};
			for (_sv2v_strm_BEEC1_idx = 0; _sv2v_strm_BEEC1_idx <= 7; _sv2v_strm_BEEC1_idx = _sv2v_strm_BEEC1_idx + 1)
				_sv2v_strm_BEEC1_out[7 - _sv2v_strm_BEEC1_idx-:1] = _sv2v_strm_BEEC1_inp[_sv2v_strm_BEEC1_idx+:1];
			_sv2v_strm_D90CD = _sv2v_strm_BEEC1_out << 0;
		end
	endfunction
	assign TransmitDataEndian = (Format[0] ? _sv2v_strm_D90CD({TransmitReadData[7:0]}) : TransmitReadData[7:0]);
	always @(posedge PCLK)
		if (~PRESETn)
			TransmitReg <= 8'b00000000;
		else if (TransmitLoad)
			TransmitReg <= TransmitDataEndian;
		else if (ShiftEdge)
			TransmitReg <= {TransmitReg[6:0], TransmitReg[0]};
	assign SPIOut = TransmitReg[7];
	assign ShiftIn = (P[2178] ? SPIOut : SPIIn);
	always @(posedge PCLK)
		if (~PRESETn)
			ReceiveShiftReg <= 8'b00000000;
		else if (SampleEdge)
			ReceiveShiftReg <= {ReceiveShiftReg[6:0], ShiftIn};
	assign LeftShiftAmount = 4'h8 - FrameLength;
	assign ASR = ReceiveShiftReg << LeftShiftAmount[2:0];
	function automatic [7:0] _sv2v_strm_A7A5E;
		input reg [7:0] inp;
		reg [7:0] _sv2v_strm_BEEC1_inp;
		reg [7:0] _sv2v_strm_BEEC1_out;
		integer _sv2v_strm_BEEC1_idx;
		begin
			_sv2v_strm_BEEC1_inp = {inp};
			for (_sv2v_strm_BEEC1_idx = 0; _sv2v_strm_BEEC1_idx <= 7; _sv2v_strm_BEEC1_idx = _sv2v_strm_BEEC1_idx + 1)
				_sv2v_strm_BEEC1_out[7 - _sv2v_strm_BEEC1_idx-:1] = _sv2v_strm_BEEC1_inp[_sv2v_strm_BEEC1_idx+:1];
			_sv2v_strm_A7A5E = _sv2v_strm_BEEC1_out << 0;
		end
	endfunction
	assign ReceiveShiftRegEndian = (Format[0] ? _sv2v_strm_A7A5E({ASR[7:0]}) : ASR[7:0]);
	assign SPIIntr = |(InterruptPending & InterruptEnable);
	assign ChipSelectInternal = (InactiveState ? ChipSelectDef : ~ChipSelectDef);
	always @(*) begin
		if (_sv2v_0)
			;
		case (ChipSelectID[1:0])
			2'b00: ChipSelectAuto = {ChipSelectDef[3], ChipSelectDef[2], ChipSelectDef[1], ChipSelectInternal[0]};
			2'b01: ChipSelectAuto = {ChipSelectDef[3], ChipSelectDef[2], ChipSelectInternal[1], ChipSelectDef[0]};
			2'b10: ChipSelectAuto = {ChipSelectDef[3], ChipSelectInternal[2], ChipSelectDef[1], ChipSelectDef[0]};
			2'b11: ChipSelectAuto = {ChipSelectInternal[3], ChipSelectDef[2], ChipSelectDef[1], ChipSelectDef[0]};
		endcase
	end
	assign SPICS = (ChipSelectMode[0] ? ChipSelectDef : ChipSelectAuto);
	initial _sv2v_0 = 0;
endmodule
module spi_controller (
	PCLK,
	PRESETn,
	TransmitStart,
	TransmitRegLoaded,
	ResetSCLKenable,
	SckDiv,
	SckMode,
	CSMode,
	Delay0,
	Delay1,
	FrameLength,
	TransmitFIFOEmpty,
	SCLKenable,
	ShiftEdge,
	SampleEdge,
	EndOfFrame,
	Transmitting,
	InactiveState,
	SPICLK
);
	reg _sv2v_0;
	input wire PCLK;
	input wire PRESETn;
	input wire TransmitStart;
	input wire TransmitRegLoaded;
	input wire ResetSCLKenable;
	input wire [11:0] SckDiv;
	input wire [1:0] SckMode;
	input wire [1:0] CSMode;
	input wire [15:0] Delay0;
	input wire [15:0] Delay1;
	input wire [3:0] FrameLength;
	input wire TransmitFIFOEmpty;
	output wire SCLKenable;
	output reg ShiftEdge;
	output reg SampleEdge;
	output reg EndOfFrame;
	output wire Transmitting;
	output wire InactiveState;
	output reg SPICLK;
	localparam HOLDMODE = 2'b10;
	localparam AUTOMODE = 2'b00;
	localparam OFFMODE = 2'b11;
	reg [2:0] CurrState;
	reg [2:0] NextState;
	reg [11:0] DivCounter;
	reg SCK;
	wire EdgePulse;
	wire ShiftEdgePulse;
	wire SampleEdgePulse;
	wire EndOfFramePulse;
	wire InvertClock;
	reg [3:0] BitNum;
	wire LastBit;
	wire ContinueTransmit;
	wire EndTransmission;
	wire NextEndDelay;
	wire CurrentEndDelay;
	wire [7:0] cssck;
	wire [7:0] sckcs;
	wire [7:0] intercs;
	wire [7:0] interxfr;
	wire Phase;
	wire HasCSSCK;
	wire HasSCKCS;
	wire HasINTERCS;
	wire HasINTERXFR;
	wire EndOfCSSCK;
	wire EndOfSCKCS;
	wire EndOfINTERCS;
	wire EndOfINTERXFR;
	wire EndOfDelay;
	reg [7:0] DelayCounter;
	wire DelayState;
	assign cssck = Delay0[7:0];
	assign sckcs = Delay0[15:8];
	assign intercs = Delay1[7:0];
	assign interxfr = Delay1[15:8];
	assign HasCSSCK = cssck > 8'b00000000;
	assign HasSCKCS = sckcs > 8'b00000000;
	assign HasINTERCS = intercs > 8'b00000000;
	assign HasINTERXFR = interxfr > 8'b00000000;
	assign EndOfCSSCK = (DelayCounter == cssck) & (CurrState == 3'd1);
	assign EndOfSCKCS = (DelayCounter == sckcs) & (CurrState == 3'd3);
	assign EndOfINTERCS = (DelayCounter == intercs) & (CurrState == 3'd5);
	assign EndOfINTERXFR = (DelayCounter == interxfr) & (CurrState == 3'd6);
	assign EndOfDelay = ((EndOfCSSCK | EndOfSCKCS) | EndOfINTERCS) | EndOfINTERXFR;
	assign SCLKenable = DivCounter == SckDiv;
	assign ContinueTransmit = ~TransmitFIFOEmpty & EndOfFrame;
	assign EndTransmission = TransmitFIFOEmpty & EndOfFrame;
	assign Phase = SckMode[0];
	always @(posedge PCLK)
		if (~PRESETn) begin
			DivCounter <= 12'b000000000000;
			SPICLK <= SckMode[1];
			SCK <= 0;
			BitNum <= 4'h0;
			DelayCounter <= 0;
		end
		else begin
			if (TransmitStart & ~DelayState)
				SCK <= 0;
			else if (SCLKenable)
				SCK <= ~SCK;
			if ((DelayState & SCK) & SCLKenable)
				DelayCounter <= DelayCounter + 8'd1;
			else if ((SCLKenable & EndOfDelay) | Transmitting)
				DelayCounter <= 8'd0;
			if (TransmitStart & ~DelayState)
				SPICLK <= SckMode[1];
			else if (SCLKenable)
				SPICLK <= ((NextState == 3'd2) & ((~Phase & Transmitting) | Phase) ? ~SPICLK : SckMode[1]);
			if ((SCLKenable | (TransmitStart & ~DelayState)) | ResetSCLKenable)
				DivCounter <= 12'b000000000000;
			else
				DivCounter <= DivCounter + 12'd1;
			if (ShiftEdge & Transmitting)
				BitNum <= BitNum + 4'd1;
			else if (EndOfFrame)
				BitNum <= 4'b0000;
		end
	assign LastBit = BitNum == (FrameLength - 4'b0001);
	assign EdgePulse = SCLKenable & Transmitting;
	assign ShiftEdgePulse = EdgePulse & ~LastBit;
	assign SampleEdgePulse = EdgePulse & (NextState == 3'd2);
	assign EndOfFramePulse = EdgePulse & LastBit;
	assign InvertClock = ^SckMode;
	always @(negedge PCLK)
		if (~PRESETn | TransmitStart) begin
			ShiftEdge <= 0;
			SampleEdge <= 0;
			EndOfFrame <= 0;
		end
		else begin
			ShiftEdge <= (InvertClock ^ SPICLK) & ShiftEdgePulse;
			SampleEdge <= (InvertClock ^ ~SPICLK) & SampleEdgePulse;
			EndOfFrame <= (InvertClock ^ SPICLK) & EndOfFramePulse;
		end
	always @(posedge PCLK)
		if (~PRESETn)
			CurrState <= 3'd0;
		else if (SCLKenable)
			CurrState <= NextState;
	always @(*) begin
		if (_sv2v_0)
			;
		case (CurrState)
			3'd0:
				if (TransmitRegLoaded) begin
					if (~HasCSSCK)
						NextState = 3'd2;
					else
						NextState = 3'd1;
				end
				else
					NextState = 3'd0;
			3'd1:
				if (EndOfCSSCK)
					NextState = 3'd2;
				else
					NextState = 3'd1;
			3'd2:
				case (CSMode)
					AUTOMODE:
						if (EndTransmission & ~HasSCKCS)
							NextState = 3'd0;
						else if (EndOfFrame & HasSCKCS)
							NextState = 3'd3;
						else if (EndOfFrame & ~HasSCKCS)
							NextState = 3'd5;
						else
							NextState = 3'd2;
					HOLDMODE:
						if (EndOfFrame & HasINTERXFR)
							NextState = 3'd6;
						else if (EndTransmission)
							NextState = 3'd4;
						else
							NextState = 3'd2;
					OFFMODE:
						if (EndOfFrame & HasINTERXFR)
							NextState = 3'd6;
						else if (EndTransmission)
							NextState = 3'd4;
						else
							NextState = 3'd2;
					default: NextState = 3'd2;
				endcase
			3'd3:
				if (EndOfSCKCS)
					NextState = 3'd5;
				else
					NextState = 3'd3;
			3'd4:
				if (CSMode == AUTOMODE)
					NextState = 3'd0;
				else if (TransmitRegLoaded)
					NextState = 3'd2;
				else
					NextState = 3'd4;
			3'd5:
				if (EndOfINTERCS) begin
					if (TransmitRegLoaded) begin
						if (HasCSSCK)
							NextState = 3'd1;
						else
							NextState = 3'd2;
					end
					else
						NextState = 3'd0;
				end
				else
					NextState = 3'd5;
			3'd6:
				if (EndOfINTERXFR) begin
					if (TransmitRegLoaded)
						NextState = 3'd2;
					else
						NextState = 3'd4;
				end
				else
					NextState = 3'd6;
			default: NextState = 3'd0;
		endcase
	end
	assign Transmitting = CurrState == 3'd2;
	assign DelayState = (((CurrState == 3'd1) | (CurrState == 3'd3)) | (CurrState == 3'd5)) | (CurrState == 3'd6);
	assign InactiveState = (CurrState == 3'd0) | (CurrState == 3'd5);
	initial _sv2v_0 = 0;
endmodule
module spi_fifo (
	PCLK,
	wen,
	ren,
	PRESETn,
	winc,
	rinc,
	wdata,
	wwatermarklevel,
	rwatermarklevel,
	rdata,
	wfull,
	rempty,
	wwatermark,
	rwatermark
);
	parameter M = 3;
	parameter N = 8;
	input wire PCLK;
	input wire wen;
	input wire ren;
	input wire PRESETn;
	input wire winc;
	input wire rinc;
	input wire [N - 1:0] wdata;
	input wire [M - 1:0] wwatermarklevel;
	input wire [M - 1:0] rwatermarklevel;
	output wire [N - 1:0] rdata;
	output reg wfull;
	output reg rempty;
	output wire wwatermark;
	output wire rwatermark;
	reg [N - 1:0] mem [0:(2 ** M) - 1];
	reg [M:0] rptr;
	reg [M:0] wptr;
	wire [M:0] rptrnext;
	wire [M:0] wptrnext;
	wire [M - 1:0] raddr;
	wire [M - 1:0] waddr;
	wire [M - 1:0] numVals;
	assign numVals = waddr - raddr;
	assign rdata = mem[raddr];
	always @(posedge PCLK)
		if ((winc & wen) & ~wfull)
			mem[waddr] <= wdata;
	always @(posedge PCLK)
		if (~PRESETn) begin
			rptr <= 1'sb0;
			wptr <= 1'sb0;
			wfull <= 1'b0;
			rempty <= 1'b1;
		end
		else begin
			if (wen) begin
				wfull <= {~wptrnext[M], wptrnext[M - 1:0]} == rptr;
				wptr <= wptrnext;
			end
			if (ren) begin
				rptr <= rptrnext;
				rempty <= wptr == rptrnext;
			end
		end
	assign raddr = rptr[M - 1:0];
	assign rptrnext = rptr + {{M {1'b0}}, rinc & ~rempty};
	assign rwatermark = ((waddr - raddr) < rwatermarklevel) & ~wfull;
	assign waddr = wptr[M - 1:0];
	assign wwatermark = ((waddr - raddr) > wwatermarklevel) | wfull;
	assign wptrnext = wptr + {{M {1'b0}}, winc & ~wfull};
endmodule
module uartPC16550D (
	PCLK,
	PRESETn,
	A,
	Din,
	Dout,
	MEMRb,
	MEMWb,
	INTR,
	TXRDYb,
	RXRDYb,
	BAUDOUTb,
	RCLK,
	SIN,
	DSRb,
	DCDb,
	CTSb,
	RIb,
	SOUT,
	RTSb,
	DTRb,
	OUT1b,
	OUT2b
);
	reg _sv2v_0;
	parameter UART_PRESCALE = 0;
	input wire PCLK;
	input wire PRESETn;
	input wire [2:0] A;
	input wire [7:0] Din;
	output reg [7:0] Dout;
	input wire MEMRb;
	input wire MEMWb;
	output reg INTR;
	output reg TXRDYb;
	output reg RXRDYb;
	output wire BAUDOUTb;
	input wire RCLK;
	input wire SIN;
	input wire DSRb;
	input wire DCDb;
	input wire CTSb;
	input wire RIb;
	output wire SOUT;
	output wire RTSb;
	output wire DTRb;
	output wire OUT1b;
	output wire OUT2b;
	localparam UART_DLL_RBR = 3'b000;
	localparam UART_DLM_IER = 3'b001;
	localparam UART_IIR = 3'b010;
	localparam UART_LCR = 3'b011;
	localparam UART_MCR = 3'b100;
	localparam UART_LSR = 3'b101;
	localparam UART_MSR = 3'b110;
	localparam UART_SCR = 3'b111;
	reg [10:0] RBR;
	reg [7:0] FCR;
	reg [7:0] LCR;
	reg [7:0] LSR;
	reg [7:0] SCR;
	reg [7:0] DLL;
	reg [7:0] DLM;
	reg [3:0] IER;
	reg [3:0] MSR;
	reg [4:0] MCR;
	reg SINd;
	reg DSRbd;
	reg DCDbd;
	reg CTSbd;
	reg RIbd;
	reg SINsync;
	reg DSRbsync;
	reg DCDbsync;
	reg CTSbsync;
	reg RIbsync;
	reg DSRb2;
	reg DCDb2;
	reg CTSb2;
	reg RIb2;
	wire SOUTbit;
	wire loop;
	wire DLAB;
	reg baudpulse;
	wire txbaudpulse;
	wire rxbaudpulse;
	reg [(16 + UART_PRESCALE) - 1:0] baudcount;
	reg [3:0] rxoversampledcnt;
	reg [3:0] txoversampledcnt;
	reg [3:0] rxbitsreceived;
	reg [3:0] txbitssent;
	reg [1:0] rxstate;
	reg [1:0] txstate;
	reg [9:0] rxshiftreg;
	reg [10:0] rxfifo [15:0];
	reg [7:0] txfifo [15:0];
	wire [4:0] rxfifotailunwrapped;
	reg [3:0] rxfifohead;
	reg [3:0] rxfifotail;
	reg [3:0] txfifohead;
	reg [3:0] txfifotail;
	reg [3:0] rxfifotriggerlevel;
	wire [3:0] rxfifoentries;
	wire [3:0] rxbitsexpected;
	wire [3:0] txbitsexpected;
	reg [10:0] RXBR;
	reg [9:0] rxtimeoutcnt;
	wire rxcentered;
	wire rxparity;
	wire rxparitybit;
	wire rxstopbit;
	wire rxparityerr;
	wire rxoverrunerr;
	wire rxframingerr;
	wire rxbreak;
	wire rxfifohaserr;
	reg rxdataready;
	wire rxfifoempty;
	wire rxfifotriggered;
	wire rxfifotimeout;
	reg rxfifodmaready;
	reg [8:0] rxdata9;
	wire [7:0] rxdata;
	wire [15:0] RXerrbit;
	wire [15:0] rxfullbit;
	wire [31:0] rxfullbitunwrapped;
	reg [7:0] TXHR;
	reg [7:0] nexttxdata;
	reg [11:0] txdata;
	reg [11:0] txsr;
	wire txnextbit;
	reg txhrfull;
	reg txsrfull;
	reg txparity;
	wire txfifoempty;
	wire txfifofull;
	reg txfifodmaready;
	wire fifoenabled;
	wire fifodmamodesel;
	wire evenparitysel;
	wire RXerr;
	wire RXerrIP;
	wire squashRXerrIP;
	wire prevSquashRXerrIP;
	wire setSquashRXerrIP;
	wire resetSquashRXerrIP;
	wire THRE;
	wire THRE_IP;
	wire squashTHRE_IP;
	wire prevSquashTHRE_IP;
	wire setSquashTHRE_IP;
	wire resetSquashTHRE_IP;
	wire rxdataavailintr;
	wire modemstatusintr;
	reg intrpending;
	reg [2:0] intrID;
	wire baudpulseComb;
	reg HeadPointerLastMove;
	always @(posedge PCLK) begin
		{SINd, DSRbd, DCDbd, CTSbd, RIbd} <= {SIN, DSRb, DCDb, CTSb, RIb};
		{SINsync, DSRbsync, DCDbsync, CTSbsync, RIbsync} <= (loop ? {SOUTbit, ~MCR[0], ~MCR[3], ~MCR[1], ~MCR[2]} : {SINd, DSRbd, DCDbd, CTSbd, RIbd});
		{DSRb2, DCDb2, CTSb2, RIb2} <= {DSRbsync, DCDbsync, CTSbsync, RIbsync};
	end
	always @(posedge PCLK)
		if (~PRESETn) begin
			IER <= 4'b0000;
			FCR <= 8'b00000000;
			LCR <= 8'b00000011;
			MCR <= 5'b00000;
			LSR <= 8'b01100000;
			MSR <= 4'b0000;
			DLL <= 8'd1;
			DLM <= 8'b00000000;
			SCR <= 8'b00000000;
		end
		else begin
			if (~MEMWb)
				case (A)
					UART_DLL_RBR:
						if (DLAB)
							DLL <= Din;
					UART_DLM_IER:
						if (DLAB)
							DLM <= Din;
						else
							IER <= Din[3:0];
					UART_IIR: FCR <= {Din[7:6], 2'b00, Din[3], 2'b00, Din[0]};
					UART_LCR: LCR <= Din;
					UART_MCR: MCR <= Din[4:0];
					UART_SCR: SCR <= Din;
				endcase
			if (~MEMWb & (A == UART_LSR))
				LSR[6:1] <= Din[6:1];
			else begin
				LSR[0] <= rxdataready;
				LSR[1] <= (LSR[1] | RXBR[10]) & ~squashRXerrIP;
				LSR[2] <= (LSR[2] | RXBR[9]) & ~squashRXerrIP;
				LSR[3] <= (LSR[3] | RXBR[8]) & ~squashRXerrIP;
				LSR[4] <= (LSR[4] | rxbreak) & ~squashRXerrIP;
				LSR[5] <= THRE;
				LSR[6] <= ~txsrfull & THRE;
				if (rxfifohaserr)
					LSR[7] <= 1'b1;
			end
			if (~MEMWb & (A == UART_MSR))
				MSR <= Din[3:0];
			else if (~MEMRb & (A == UART_MSR))
				MSR <= 4'b0000;
			else begin
				MSR[0] <= MSR[0] | (CTSb2 ^ CTSbsync);
				MSR[1] <= MSR[1] | (DSRb2 ^ DSRbsync);
				MSR[2] <= MSR[2] | (~RIb2 & RIbsync);
				MSR[3] <= MSR[3] | (DCDb2 ^ DCDbsync);
			end
		end
	always @(*) begin
		if (_sv2v_0)
			;
		if (~MEMRb)
			case (A)
				UART_DLL_RBR:
					if (DLAB)
						Dout = DLL;
					else
						Dout = RBR[7:0];
				UART_DLM_IER:
					if (DLAB)
						Dout = DLM;
					else
						Dout = {4'b0000, IER[3:0]};
				UART_IIR: Dout = {{2 {fifoenabled}}, 2'b00, intrID[2:0], ~intrpending};
				UART_LCR: Dout = LCR;
				UART_MCR: Dout = {3'b000, MCR};
				UART_LSR: Dout = LSR;
				UART_MSR: Dout = {~DCDbsync, ~RIbsync, ~DSRbsync, ~CTSbsync, MSR[3:0]};
				UART_SCR: Dout = SCR;
			endcase
		else
			Dout = 8'b00000000;
	end
	always @(posedge PCLK)
		if (~PRESETn) begin
			baudcount <= 1;
			baudpulse <= 1'b0;
		end
		else if ((~MEMWb & DLAB) & ((A == 3'b000) | (A == 3'b001)))
			baudcount <= 1;
		else begin
			baudpulse <= baudpulseComb;
			baudcount <= (baudpulseComb ? 1 : baudcount + 1);
		end
	assign baudpulseComb = baudcount == {DLM, DLL, {UART_PRESCALE {1'b0}}};
	assign txbaudpulse = baudpulse;
	assign BAUDOUTb = ~baudpulse;
	assign rxbaudpulse = ~RCLK;
	always @(posedge PCLK)
		if (~PRESETn) begin
			rxoversampledcnt <= 1'sb0;
			rxstate <= 2'd0;
			rxbitsreceived <= 1'sb0;
			rxtimeoutcnt <= 1'sb0;
		end
		else begin
			if ((rxstate == 2'd0) & ~SINsync) begin
				rxstate <= 2'd1;
				rxoversampledcnt <= 1'sb0;
				rxbitsreceived <= 1'sb0;
				if (~rxfifotimeout)
					rxtimeoutcnt <= 1'sb0;
			end
			else if (rxbaudpulse & (rxstate == 2'd1)) begin
				rxoversampledcnt <= rxoversampledcnt + 4'b0001;
				if (rxcentered)
					rxbitsreceived <= rxbitsreceived + 1;
				if (rxbitsreceived == rxbitsexpected)
					rxstate <= 2'd2;
			end
			else if ((rxstate == 2'd2) | (rxstate == 2'd3)) begin
				if (rxbreak & ~SINsync)
					rxstate <= 2'd3;
				else
					rxstate <= 2'd0;
			end
			if ((~MEMRb & (A == 3'b000)) & ~DLAB)
				rxtimeoutcnt <= 1'sb0;
			else if (((fifoenabled & ~rxfifoempty) & rxbaudpulse) & ~rxfifotimeout)
				rxtimeoutcnt <= rxtimeoutcnt + 1;
		end
	assign rxcentered = rxbaudpulse & (rxoversampledcnt == 4'b1000);
	assign rxbitsexpected = (((4'd1 + 4'd5) + {2'b00, LCR[1:0]}) + {3'b000, LCR[3]}) + 4'd1;
	always @(posedge PCLK)
		if (~PRESETn)
			rxshiftreg <= 10'b0000000001;
		else if (rxcentered)
			rxshiftreg <= {rxshiftreg[8:0], SINsync};
	assign rxparitybit = rxshiftreg[1];
	assign rxstopbit = rxshiftreg[0];
	always @(*) begin
		if (_sv2v_0)
			;
		case (LCR[1:0])
			2'b00: rxdata9 = {3'b000, rxshiftreg[1], rxshiftreg[2], rxshiftreg[3], rxshiftreg[4], rxshiftreg[5], rxshiftreg[6]};
			2'b01: rxdata9 = {2'b00, rxshiftreg[1], rxshiftreg[2], rxshiftreg[3], rxshiftreg[4], rxshiftreg[5], rxshiftreg[6], rxshiftreg[7]};
			2'b10: rxdata9 = {1'b0, rxshiftreg[1], rxshiftreg[2], rxshiftreg[3], rxshiftreg[4], rxshiftreg[5], rxshiftreg[6], rxshiftreg[7], rxshiftreg[8]};
			2'b11: rxdata9 = {rxshiftreg[1], rxshiftreg[2], rxshiftreg[3], rxshiftreg[4], rxshiftreg[5], rxshiftreg[6], rxshiftreg[7], rxshiftreg[8], rxshiftreg[9]};
		endcase
	end
	assign rxdata = (LCR[3] ? rxdata9[7:0] : rxdata9[8:1]);
	assign rxparity = ^rxdata;
	assign rxparityerr = ((rxparity ^ rxparitybit) ^ ~evenparitysel) & LCR[3];
	assign rxoverrunerr = (fifoenabled ? rxfifoentries == 15 : rxdataready);
	assign rxframingerr = ~rxstopbit;
	assign rxbreak = rxframingerr & (rxdata9 == 9'b000000000);
	always @(posedge PCLK)
		if (~PRESETn) begin
			rxfifohead <= 1'sb0;
			rxfifotail <= 1'sb0;
			rxdataready <= 1'b0;
			RXBR <= 1'sb0;
		end
		else if ((~MEMWb & (A == 3'b010)) & Din[1]) begin
			rxfifohead <= 1'sb0;
			rxfifotail <= 1'sb0;
			rxdataready <= 1'b0;
		end
		else if (rxstate == 2'd2) begin
			RXBR <= {rxoverrunerr, rxparityerr, rxframingerr, rxdata};
			if (fifoenabled) begin
				rxfifo[rxfifohead] <= {rxoverrunerr, rxparityerr, rxframingerr, rxdata};
				rxfifohead <= rxfifohead + 1'b1;
			end
			rxdataready <= 1'b1;
		end
		else if ((~MEMRb & (A == 3'b000)) & ~DLAB) begin
			if (fifoenabled) begin
				if (~rxfifoempty)
					rxfifotail <= rxfifotail + 1;
				if (rxfifoentries == 1)
					rxdataready <= 1'b0;
			end
			else begin
				rxdataready <= 1'b0;
				RXBR <= {1'b0, RXBR[9:0]};
			end
		end
		else if (~MEMWb & (A == 3'b010)) begin
			if (Din[1] | ~Din[0]) begin
				rxfifohead <= 1'sb0;
				rxfifotail <= 1'sb0;
			end
		end
	assign rxfifoempty = rxfifohead == rxfifotail;
	assign rxfifoentries = (rxfifohead >= rxfifotail ? rxfifohead - rxfifotail : (rxfifohead + 16) - rxfifotail);
	assign rxfifotriggered = rxfifoentries >= rxfifotriggerlevel;
	assign rxfifotimeout = rxtimeoutcnt == {rxbitsexpected, 6'b000000};
	assign rxfifotailunwrapped = (rxfifotail < rxfifohead ? {1'b1, rxfifotail} : {1'b0, rxfifotail});
	genvar _gv_i_6;
	generate
		for (_gv_i_6 = 0; _gv_i_6 < 32; _gv_i_6 = _gv_i_6 + 1) begin : rxfull
			localparam i = _gv_i_6;
			if (i == 0) begin : genblk1
				assign rxfullbitunwrapped[i] = (rxfifohead == 0) & (rxfifotail != 0);
			end
			else begin : genblk1
				assign rxfullbitunwrapped[i] = (({1'b0, rxfifohead} == i) | rxfullbitunwrapped[i - 1]) & (rxfifotailunwrapped != i);
			end
		end
		for (_gv_i_6 = 0; _gv_i_6 < 16; _gv_i_6 = _gv_i_6 + 1) begin : rx
			localparam i = _gv_i_6;
			assign RXerrbit[i] = |rxfifo[i][10:8];
			assign rxfullbit[i] = rxfullbitunwrapped[i] | rxfullbitunwrapped[i + 16];
		end
	endgenerate
	assign rxfifohaserr = |(RXerrbit & rxfullbit);
	always @(posedge PCLK)
		if (~PRESETn)
			rxfifodmaready <= 1'b0;
		else if (rxfifotriggered | rxfifotimeout)
			rxfifodmaready <= 1'b1;
		else if (rxfifoempty)
			rxfifodmaready <= 1'b0;
	always @(*) begin
		if (_sv2v_0)
			;
		if (fifoenabled) begin
			if (rxfifoempty)
				RBR = 11'b00000000000;
			else
				RBR = rxfifo[rxfifotail];
			if (fifodmamodesel)
				RXRDYb = ~rxfifodmaready;
			else
				RXRDYb = rxfifoempty;
		end
		else begin
			RBR = RXBR;
			RXRDYb = ~rxdataready;
		end
	end
	always @(posedge PCLK)
		if (~PRESETn) begin
			txoversampledcnt <= 1'sb0;
			txstate <= 2'd0;
			txbitssent <= 1'sb0;
		end
		else if ((txstate == 2'd0) & txsrfull) begin
			txstate <= 2'd1;
			txoversampledcnt <= 4'b0001;
			txbitssent <= 1'sb0;
		end
		else if (txbaudpulse & (txstate == 2'd1)) begin
			txoversampledcnt <= txoversampledcnt + 1'b1;
			if (txnextbit) begin
				txbitssent <= txbitssent + 1'b1;
				if (txbitssent == txbitsexpected)
					txstate <= 2'd2;
			end
		end
		else if (txstate == 2'd2)
			txstate <= 2'd0;
	assign txbitsexpected = (((((4'd1 + 4'd5) + {2'b00, LCR[1:0]}) + {3'b000, LCR[3]}) + 4'd1) + {3'b000, LCR[2]}) - 4'd1;
	assign txnextbit = txbaudpulse & (txoversampledcnt == 4'b0000);
	always @(*) begin
		if (_sv2v_0)
			;
		nexttxdata = (fifoenabled ? txfifo[txfifotail] : TXHR);
		case (LCR[1:0])
			2'b00: txparity = ^nexttxdata[4:0] ^ ~evenparitysel;
			2'b01: txparity = ^nexttxdata[5:0] ^ ~evenparitysel;
			2'b10: txparity = ^nexttxdata[6:0] ^ ~evenparitysel;
			2'b11: txparity = ^nexttxdata[7:0] ^ ~evenparitysel;
		endcase
		case ({LCR[3], LCR[1:0]})
			3'b000: txdata = {1'b0, nexttxdata[0], nexttxdata[1], nexttxdata[2], nexttxdata[3], nexttxdata[4], 6'b111111};
			3'b001: txdata = {1'b0, nexttxdata[0], nexttxdata[1], nexttxdata[2], nexttxdata[3], nexttxdata[4], nexttxdata[5], 5'b11111};
			3'b010: txdata = {1'b0, nexttxdata[0], nexttxdata[1], nexttxdata[2], nexttxdata[3], nexttxdata[4], nexttxdata[5], nexttxdata[6], 4'b1111};
			3'b011: txdata = {1'b0, nexttxdata[0], nexttxdata[1], nexttxdata[2], nexttxdata[3], nexttxdata[4], nexttxdata[5], nexttxdata[6], nexttxdata[7], 3'b111};
			3'b100: txdata = {1'b0, nexttxdata[0], nexttxdata[1], nexttxdata[2], nexttxdata[3], nexttxdata[4], txparity, 5'b11111};
			3'b101: txdata = {1'b0, nexttxdata[0], nexttxdata[1], nexttxdata[2], nexttxdata[3], nexttxdata[4], nexttxdata[5], txparity, 4'b1111};
			3'b110: txdata = {1'b0, nexttxdata[0], nexttxdata[1], nexttxdata[2], nexttxdata[3], nexttxdata[4], nexttxdata[5], nexttxdata[6], txparity, 3'b111};
			3'b111: txdata = {1'b0, nexttxdata[0], nexttxdata[1], nexttxdata[2], nexttxdata[3], nexttxdata[4], nexttxdata[5], nexttxdata[6], nexttxdata[7], txparity, 2'b11};
		endcase
	end
	always @(posedge PCLK)
		if (~PRESETn) begin
			txfifohead <= 1'sb0;
			txfifotail <= 1'sb0;
			txhrfull <= 1'b0;
			txsrfull <= 1'b0;
			TXHR <= 1'sb0;
			txsr <= 12'hfff;
		end
		else if ((~MEMWb & (A == 3'b010)) & Din[2]) begin
			txfifohead <= 1'sb0;
			txfifotail <= 1'sb0;
		end
		else begin
			if ((~MEMWb & (A == 3'b000)) & ~DLAB) begin
				if (fifoenabled) begin
					txfifo[txfifohead] <= Din;
					txfifohead <= txfifohead + 4'b0001;
				end
				else begin
					TXHR <= Din;
					txhrfull <= 1'b1;
				end
				$write("%c", Din);
			end
			if (txstate == 2'd0) begin
				if (fifoenabled) begin
					if (~txfifoempty & ~txsrfull) begin
						txsr <= txdata;
						txfifotail <= txfifotail + 1;
						txsrfull <= 1'b1;
					end
				end
				else if (txhrfull) begin
					txsr <= txdata;
					txhrfull <= 1'b0;
					txsrfull <= 1'b1;
				end
			end
			else if (txstate == 2'd2)
				txsrfull <= 1'b0;
			else if ((txstate == 2'd1) & txnextbit)
				txsr <= {txsr[10:0], 1'b1};
			if (!MEMWb & (A == 3'b010)) begin
				if (Din[2] | ~Din[0]) begin
					txfifohead <= 1'sb0;
					txfifotail <= 1'sb0;
				end
			end
		end
	always @(posedge PCLK)
		if (~PRESETn)
			HeadPointerLastMove <= 1'b0;
		else if (((fifoenabled & ~MEMWb) & (A == 3'b000)) & ~DLAB)
			HeadPointerLastMove <= 1'b1;
		else if (((fifoenabled & ~txfifoempty) & ~txsrfull) & (txstate == 2'd0))
			HeadPointerLastMove <= 1'b0;
	assign txfifoempty = (txfifohead == txfifotail) & ~HeadPointerLastMove;
	assign txfifofull = (txfifohead == txfifotail) & HeadPointerLastMove;
	always @(posedge PCLK)
		if (~PRESETn)
			txfifodmaready <= 1'b0;
		else if (txfifoempty)
			txfifodmaready <= 1'b1;
		else if (txfifofull)
			txfifodmaready <= 1'b0;
	always @(*) begin
		if (_sv2v_0)
			;
		if (fifoenabled & fifodmamodesel)
			TXRDYb = ~txfifodmaready;
		else
			TXRDYb = ~THRE;
	end
	assign SOUTbit = txsr[11];
	assign SOUT = (loop ? 1 : (LCR[6] ? 1'b0 : SOUTbit));
	assign RXerr = |LSR[4:1];
	assign RXerrIP = RXerr & ~squashRXerrIP;
	assign rxdataavailintr = (fifoenabled ? rxfifotriggered : rxdataready);
	assign THRE = (fifoenabled ? txfifoempty : ~txhrfull);
	assign THRE_IP = THRE & ~squashTHRE_IP;
	assign modemstatusintr = |MSR[3:0];
	always @(*) begin
		if (_sv2v_0)
			;
		intrpending = 1'b1;
		if (RXerrIP & IER[2])
			intrID = 3'b011;
		else if (rxdataavailintr & IER[0])
			intrID = 3'b010;
		else if ((rxfifotimeout & fifoenabled) & IER[0])
			intrID = 3'b110;
		else if (THRE_IP & IER[1])
			intrID = 3'b001;
		else if (modemstatusintr & IER[3])
			intrID = 3'b000;
		else begin
			intrID = 3'b000;
			intrpending = 1'b0;
		end
	end
	always @(posedge PCLK) INTR <= intrpending;
	assign setSquashRXerrIP = ~MEMRb & (A == 3'b101);
	assign resetSquashRXerrIP = rxstate == 2'd2;
	assign squashRXerrIP = (prevSquashRXerrIP | setSquashRXerrIP) & ~resetSquashRXerrIP;
	flopr #(.WIDTH(1)) squashRXerrIPreg(
		.clk(PCLK),
		.reset(~PRESETn),
		.d(squashRXerrIP),
		.q(prevSquashRXerrIP)
	);
	assign setSquashTHRE_IP = (~MEMRb & (A == 3'b010)) & (intrID == 3'h1);
	assign resetSquashTHRE_IP = ~THRE;
	assign squashTHRE_IP = prevSquashTHRE_IP & ~resetSquashTHRE_IP;
	flopr #(.WIDTH(1)) squashTHRE_IPreg(
		.clk(PCLK),
		.reset(~PRESETn),
		.d(squashTHRE_IP | setSquashTHRE_IP),
		.q(prevSquashTHRE_IP)
	);
	assign loop = MCR[4];
	assign DTRb = ~MCR[0] | loop;
	assign RTSb = ~MCR[1] | loop;
	assign OUT1b = ~MCR[2] | loop;
	assign OUT2b = ~MCR[3] | loop;
	assign DLAB = LCR[7];
	assign evenparitysel = LCR[4];
	assign fifoenabled = FCR[0];
	assign fifodmamodesel = FCR[3];
	always @(*) begin
		if (_sv2v_0)
			;
		case (FCR[7:6])
			2'b00: rxfifotriggerlevel = 4'd1;
			2'b01: rxfifotriggerlevel = 4'd4;
			2'b10: rxfifotriggerlevel = 4'd8;
			2'b11: rxfifotriggerlevel = 4'd14;
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
module uart_apb (
	PCLK,
	PRESETn,
	PSEL,
	PADDR,
	PWDATA,
	PSTRB,
	PWRITE,
	PENABLE,
	PRDATA,
	PREADY,
	SIN,
	DSRb,
	DCDb,
	CTSb,
	RIb,
	SOUT,
	RTSb,
	DTRb,
	OUT1b,
	OUT2b,
	INTR,
	TXRDYb,
	RXRDYb
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire PCLK;
	input wire PRESETn;
	input wire PSEL;
	input wire [2:0] PADDR;
	input wire [$signed(P[4216-:32]) - 1:0] PWDATA;
	input wire [($signed(P[4216-:32]) / 8) - 1:0] PSTRB;
	input wire PWRITE;
	input wire PENABLE;
	output wire [$signed(P[4216-:32]) - 1:0] PRDATA;
	output wire PREADY;
	input wire SIN;
	input wire DSRb;
	input wire DCDb;
	input wire CTSb;
	input wire RIb;
	output wire SOUT;
	output wire RTSb;
	output wire DTRb;
	output wire OUT1b;
	output wire OUT2b;
	output wire INTR;
	output wire TXRDYb;
	output wire RXRDYb;
	wire [2:0] entry;
	wire MEMRb;
	wire MEMWb;
	wire memread;
	wire memwrite;
	wire [7:0] Din;
	wire [7:0] Dout;
	assign memwrite = (PWRITE & PENABLE) & PSEL;
	assign memread = (~PWRITE & PENABLE) & PSEL;
	assign PREADY = 1'b1;
	assign entry = PADDR[2:0];
	assign MEMRb = ~memread;
	assign MEMWb = ~memwrite;
	assign Din = PWDATA[7:0];
	generate
		if ($signed(P[4216-:32]) == 64) begin : genblk1
			assign PRDATA = {Dout, Dout, Dout, Dout, Dout, Dout, Dout, Dout};
		end
		else begin : genblk1
			assign PRDATA = {Dout, Dout, Dout, Dout};
		end
	endgenerate
	wire BAUDOUTb;
	uartPC16550D #(.UART_PRESCALE($signed(P[2177-:32]))) uartPC(
		.PCLK(PCLK),
		.PRESETn(PRESETn),
		.A(entry),
		.Din(Din),
		.Dout(Dout),
		.MEMRb(MEMRb),
		.MEMWb(MEMWb),
		.INTR(INTR),
		.TXRDYb(TXRDYb),
		.RXRDYb(RXRDYb),
		.BAUDOUTb(BAUDOUTb),
		.RCLK(BAUDOUTb),
		.SIN(SIN),
		.DSRb(DSRb),
		.DCDb(DCDb),
		.CTSb(CTSb),
		.RIb(RIb),
		.SOUT(SOUT),
		.RTSb(RTSb),
		.DTRb(DTRb),
		.OUT1b(OUT1b),
		.OUT2b(OUT2b)
	);
endmodule
module uncore (
	HCLK,
	HRESETn,
	TIMECLK,
	HADDR,
	HWDATA,
	HWSTRB,
	HWRITE,
	HSIZE,
	HBURST,
	HPROT,
	HTRANS,
	HMASTLOCK,
	HRDATAEXT,
	HREADYEXT,
	HRESPEXT,
	HRDATA,
	HREADY,
	HRESP,
	HSELEXT,
	MTimerInt,
	MSwInt,
	MExtInt,
	SExtInt,
	MTIME_CLINT,
	GPIOIN,
	GPIOOUT,
	GPIOEN,
	UARTSin,
	UARTSout,
	SPIIn,
	SPIOut,
	SPICS,
	SPICLK,
	SDCIn,
	SDCCmd,
	SDCCS,
	SDCCLK
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire HCLK;
	input wire HRESETn;
	input wire TIMECLK;
	input wire [$signed(P[1640-:32]) - 1:0] HADDR;
	input wire [$signed(P[4151-:32]) - 1:0] HWDATA;
	input wire [($signed(P[4216-:32]) / 8) - 1:0] HWSTRB;
	input wire HWRITE;
	input wire [2:0] HSIZE;
	input wire [2:0] HBURST;
	input wire [3:0] HPROT;
	input wire [1:0] HTRANS;
	input wire HMASTLOCK;
	input wire [$signed(P[4151-:32]) - 1:0] HRDATAEXT;
	input wire HREADYEXT;
	input wire HRESPEXT;
	output wire [$signed(P[4151-:32]) - 1:0] HRDATA;
	output wire HREADY;
	output wire HRESP;
	output wire HSELEXT;
	output wire MTimerInt;
	output wire MSwInt;
	output wire MExtInt;
	output wire SExtInt;
	output wire [63:0] MTIME_CLINT;
	input wire [31:0] GPIOIN;
	output wire [31:0] GPIOOUT;
	output wire [31:0] GPIOEN;
	input wire UARTSin;
	output wire UARTSout;
	input wire SPIIn;
	output wire SPIOut;
	output wire [3:0] SPICS;
	output wire SPICLK;
	input wire SDCIn;
	output wire SDCCmd;
	output wire [3:0] SDCCS;
	output wire SDCCLK;
	wire [$signed(P[4216-:32]) - 1:0] HREADRam;
	wire [$signed(P[4216-:32]) - 1:0] HREADSDC;
	wire [11:0] HSELRegions;
	wire HSELDTIM;
	wire HSELIROM;
	wire HSELRam;
	wire HSELCLINT;
	wire HSELPLIC;
	wire HSELGPIO;
	wire HSELUART;
	wire HSELSDC;
	wire HSELSPI;
	wire HSELDTIMD;
	wire HSELIROMD;
	wire HSELEXTD;
	wire HSELRamD;
	wire HSELCLINTD;
	wire HSELPLICD;
	wire HSELGPIOD;
	wire HSELUARTD;
	wire HSELSDCD;
	wire HSELSPID;
	wire HRESPRam;
	wire HRESPSDC;
	wire HREADYRam;
	wire HRESPSDCD;
	wire [$signed(P[4216-:32]) - 1:0] HREADBootRom;
	wire HSELBootRom;
	wire HSELBootRomD;
	wire HRESPBootRom;
	wire HREADYBootRom;
	wire HREADYSDC;
	wire HSELNoneD;
	wire UARTIntr;
	wire GPIOIntr;
	wire SPIIntr;
	wire SDCIntM;
	wire PCLK;
	wire PRESETn;
	wire PWRITE;
	wire PENABLE;
	wire [5:0] PSEL;
	wire [31:0] PADDR;
	wire [$signed(P[4216-:32]) - 1:0] PWDATA;
	wire [($signed(P[4216-:32]) / 8) - 1:0] PSTRB;
	wire [5:0] PREADY;
	wire [(6 * $signed(P[4216-:32])) - 1:0] PRDATA;
	wire [$signed(P[4216-:32]) - 1:0] HREADBRIDGE;
	wire HRESPBRIDGE;
	wire HREADYBRIDGE;
	wire HSELBRIDGE;
	wire HSELBRIDGED;
	wire SDCIntr;
	adrdecs #(.P(P)) adrdecs(
		.PhysicalAddress(HADDR),
		.AccessRW(1'b1),
		.AccessRX(1'b1),
		.AccessRWXC(1'b1),
		.Size(HSIZE[1:0]),
		.SelRegions(HSELRegions)
	);
	assign {HSELSPI, HSELSDC, HSELPLIC, HSELUART, HSELGPIO, HSELCLINT, HSELRam, HSELBootRom, HSELEXT, HSELIROM, HSELDTIM} = HSELRegions[11:1];
	ahbapbbridge #(
		.P(P),
		.PERIPHS(6)
	) ahbapbbridge(
		.HCLK(HCLK),
		.HRESETn(HRESETn),
		.HSEL({HSELSDC, HSELSPI, HSELUART, HSELPLIC, HSELCLINT, HSELGPIO}),
		.HADDR(HADDR),
		.HWDATA(HWDATA),
		.HWSTRB(HWSTRB),
		.HWRITE(HWRITE),
		.HTRANS(HTRANS),
		.HREADY(HREADY),
		.HRDATA(HREADBRIDGE),
		.HRESP(HRESPBRIDGE),
		.HREADYOUT(HREADYBRIDGE),
		.PCLK(PCLK),
		.PRESETn(PRESETn),
		.PSEL(PSEL),
		.PWRITE(PWRITE),
		.PENABLE(PENABLE),
		.PADDR(PADDR),
		.PWDATA(PWDATA),
		.PSTRB(PSTRB),
		.PREADY(PREADY),
		.PRDATA(PRDATA)
	);
	assign HSELBRIDGE = ((((HSELGPIO | HSELCLINT) | HSELPLIC) | HSELUART) | HSELSPI) | HSELSDC;
	generate
		if (P[3212]) begin : ram
			ram_ahb #(
				.P(P),
				.RANGE(P[3147-:64]),
				.PRELOAD(P[3083])
			) ram(
				.HCLK(HCLK),
				.HRESETn(HRESETn),
				.HSELRam(HSELRam),
				.HADDR(HADDR),
				.HWRITE(HWRITE),
				.HREADY(HREADY),
				.HTRANS(HTRANS),
				.HWDATA(HWDATA),
				.HWSTRB(HWSTRB),
				.HREADRam(HREADRam),
				.HRESPRam(HRESPRam),
				.HREADYRam(HREADYRam)
			);
		end
		else begin : genblk1
			assign {HREADRam, HRESPRam, HREADYRam} = 1'sb0;
		end
		if (P[3342]) begin : bootrom
			rom_ahb #(
				.P(P),
				.RANGE(P[3277-:64]),
				.PRELOAD(P[3213])
			) bootrom(
				.HCLK(HCLK),
				.HRESETn(HRESETn),
				.HSELRom(HSELBootRom),
				.HADDR(HADDR),
				.HREADY(HREADY),
				.HTRANS(HTRANS),
				.HREADRom(HREADBootRom),
				.HRESPRom(HRESPBootRom),
				.HREADYRom(HREADYBootRom)
			);
		end
		else begin : genblk2
			assign {HREADBootRom, HRESPBootRom, HREADYBootRom} = 1'sb0;
		end
		if (P[2953] == 1) begin : clint
			clint_apb #(.P(P)) clint(
				.PCLK(PCLK),
				.PRESETn(PRESETn),
				.PSEL(PSEL[1]),
				.PADDR(PADDR[15:0]),
				.PWDATA(PWDATA),
				.PSTRB(PSTRB),
				.PWRITE(PWRITE),
				.PENABLE(PENABLE),
				.PRDATA(PRDATA[$signed(P[4216-:32])+:$signed(P[4216-:32])]),
				.PREADY(PREADY[1]),
				.MTIME(MTIME_CLINT),
				.MTimerInt(MTimerInt),
				.MSwInt(MSwInt)
			);
		end
		else begin : clint
			assign MTIME_CLINT = 1'sb0;
			assign MTimerInt = 1'b0;
			assign MSwInt = 1'b0;
		end
		if (P[2566] == 1) begin : plic
			plic_apb #(.P(P)) plic(
				.PCLK(PCLK),
				.PRESETn(PRESETn),
				.PSEL(PSEL[2]),
				.PADDR(PADDR[27:0]),
				.PWDATA(PWDATA),
				.PSTRB(PSTRB),
				.PWRITE(PWRITE),
				.PENABLE(PENABLE),
				.PRDATA(PRDATA[2 * $signed(P[4216-:32])+:$signed(P[4216-:32])]),
				.PREADY(PREADY[2]),
				.UARTIntr(UARTIntr),
				.GPIOIntr(GPIOIntr),
				.SDCIntr(SDCIntr),
				.SPIIntr(SPIIntr),
				.MExtInt(MExtInt),
				.SExtInt(SExtInt)
			);
		end
		else begin : plic
			assign MExtInt = 1'b0;
			assign SExtInt = 1'b0;
		end
		if (P[2824] == 1) begin : gpio
			gpio_apb #(.P(P)) gpio(
				.PCLK(PCLK),
				.PRESETn(PRESETn),
				.PSEL(PSEL[0]),
				.PADDR(PADDR[7:0]),
				.PWDATA(PWDATA),
				.PSTRB(PSTRB),
				.PWRITE(PWRITE),
				.PENABLE(PENABLE),
				.PRDATA(PRDATA[0+:$signed(P[4216-:32])]),
				.PREADY(PREADY[0]),
				.iof0(),
				.iof1(),
				.GPIOIN(GPIOIN),
				.GPIOOUT(GPIOOUT),
				.GPIOEN(GPIOEN),
				.GPIOIntr(GPIOIntr)
			);
		end
		else begin : gpio
			assign GPIOOUT = 1'sb0;
			assign GPIOEN = 1'sb0;
			assign GPIOIntr = 1'b0;
		end
		if (P[2695] == 1) begin : uartgen
			uart_apb #(.P(P)) uart(
				.PCLK(PCLK),
				.PRESETn(PRESETn),
				.PSEL(PSEL[3]),
				.PADDR(PADDR[2:0]),
				.PWDATA(PWDATA),
				.PSTRB(PSTRB),
				.PWRITE(PWRITE),
				.PENABLE(PENABLE),
				.PRDATA(PRDATA[3 * $signed(P[4216-:32])+:$signed(P[4216-:32])]),
				.PREADY(PREADY[3]),
				.SIN(UARTSin),
				.DSRb(1'b1),
				.DCDb(1'b1),
				.CTSb(1'b0),
				.RIb(1'b1),
				.SOUT(UARTSout),
				.RTSb(),
				.DTRb(),
				.OUT1b(),
				.OUT2b(),
				.INTR(UARTIntr),
				.TXRDYb(),
				.RXRDYb()
			);
		end
		else begin : uart
			assign UARTSout = 1'b0;
			assign UARTIntr = 1'b0;
		end
		if (P[2308] == 1) begin : spi
			spi_apb #(.P(P)) spi(
				.PCLK(PCLK),
				.PRESETn(PRESETn),
				.PSEL(PSEL[4]),
				.PADDR(PADDR[7:0]),
				.PWDATA(PWDATA),
				.PSTRB(PSTRB),
				.PWRITE(PWRITE),
				.PENABLE(PENABLE),
				.PREADY(PREADY[4]),
				.PRDATA(PRDATA[4 * $signed(P[4216-:32])+:$signed(P[4216-:32])]),
				.SPIOut(SPIOut),
				.SPIIn(SPIIn),
				.SPICS(SPICS),
				.SPICLK(SPICLK),
				.SPIIntr(SPIIntr)
			);
		end
		else begin : spi
			assign SPIOut = 1'b0;
			assign SPICS = 1'sb0;
			assign SPIIntr = 1'b0;
			assign SPICLK = 1'b0;
		end
		if (P[2437] == 1) begin : sdc
			spi_apb #(.P(P)) sdc(
				.PCLK(PCLK),
				.PRESETn(PRESETn),
				.PSEL(PSEL[5]),
				.PADDR(PADDR[7:0]),
				.PWDATA(PWDATA),
				.PSTRB(PSTRB),
				.PWRITE(PWRITE),
				.PENABLE(PENABLE),
				.PREADY(PREADY[5]),
				.PRDATA(PRDATA[5 * $signed(P[4216-:32])+:$signed(P[4216-:32])]),
				.SPIOut(SDCCmd),
				.SPIIn(SDCIn),
				.SPICS(SDCCS),
				.SPICLK(SDCCLK),
				.SPIIntr(SDCIntr)
			);
		end
		else begin : sdc
			assign SDCCmd = 1'sb0;
			assign SDCCS = 4'b0000;
			assign SDCIntr = 1'b0;
			assign SDCCLK = 1'b0;
		end
	endgenerate
	assign HRDATA = ((({$signed(P[4216-:32]) {HSELRamD}} & HREADRam) | ({$signed(P[4216-:32]) {HSELEXTD}} & HRDATAEXT)) | ({$signed(P[4216-:32]) {HSELBRIDGED}} & HREADBRIDGE)) | ({$signed(P[4216-:32]) {HSELBootRomD}} & HREADBootRom);
	assign HRESP = (((HSELRamD & HRESPRam) | (HSELEXTD & HRESPEXT)) | (HSELBRIDGE & HRESPBRIDGE)) | (HSELBootRomD & HRESPBootRom);
	assign HREADY = ((((HSELRamD & HREADYRam) | (HSELEXTD & HREADYEXT)) | (HSELBRIDGED & HREADYBRIDGE)) | (HSELBootRomD & HREADYBootRom)) | HSELNoneD;
	flopenl #(.WIDTH(12)) hseldelayreg(
		.clk(HCLK),
		.load(~HRESETn),
		.en(HREADY),
		.d(HSELRegions),
		.val(12'b000000000001),
		.q({HSELSPID, HSELSDCD, HSELPLICD, HSELUARTD, HSELGPIOD, HSELCLINTD, HSELRamD, HSELBootRomD, HSELEXTD, HSELIROMD, HSELDTIMD, HSELNoneD})
	);
	flopenr #(.WIDTH(1)) hselbridgedelayreg(
		.clk(HCLK),
		.reset(~HRESETn),
		.en(HREADY),
		.d(HSELBRIDGE),
		.q(HSELBRIDGED)
	);
endmodule
module wallypipelinedcore (
	clk,
	reset,
	MTimerInt,
	MExtInt,
	SExtInt,
	MSwInt,
	MTIME_CLINT,
	HRDATA,
	HREADY,
	HRESP,
	HCLK,
	HRESETn,
	HADDR,
	HWDATA,
	HWSTRB,
	HWRITE,
	HSIZE,
	HBURST,
	HPROT,
	HTRANS,
	HMASTLOCK,
	ExternalStall
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire MTimerInt;
	input wire MExtInt;
	input wire SExtInt;
	input wire MSwInt;
	input wire [63:0] MTIME_CLINT;
	input wire [$signed(P[4151-:32]) - 1:0] HRDATA;
	input wire HREADY;
	input wire HRESP;
	output wire HCLK;
	output wire HRESETn;
	output wire [$signed(P[1640-:32]) - 1:0] HADDR;
	output wire [$signed(P[4151-:32]) - 1:0] HWDATA;
	output wire [($signed(P[4216-:32]) / 8) - 1:0] HWSTRB;
	output wire HWRITE;
	output wire [2:0] HSIZE;
	output wire [2:0] HBURST;
	output wire [3:0] HPROT;
	output wire [1:0] HTRANS;
	output wire HMASTLOCK;
	input wire ExternalStall;
	wire StallF;
	wire StallD;
	wire StallE;
	wire StallM;
	wire StallW;
	wire FlushD;
	wire FlushE;
	wire FlushM;
	wire FlushW;
	wire TrapM;
	wire RetM;
	wire IntDivE;
	wire W64E;
	wire CSRReadM;
	wire CSRWriteM;
	wire PrivilegedM;
	wire [1:0] AtomicM;
	wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcAE;
	wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcBE;
	wire [$signed(P[4216-:32]) - 1:0] SrcAM;
	wire [2:0] Funct3E;
	wire [31:0] InstrD;
	wire [31:0] InstrM;
	wire [31:0] InstrOrigM;
	wire [$signed(P[4216-:32]) - 1:0] PCSpillF;
	wire [$signed(P[4216-:32]) - 1:0] PCE;
	wire [$signed(P[4216-:32]) - 1:0] PCLinkE;
	wire [$signed(P[4216-:32]) - 1:0] PCM;
	wire [$signed(P[4216-:32]) - 1:0] CSRReadValW;
	wire [$signed(P[4216-:32]) - 1:0] MDUResultW;
	wire [$signed(P[4216-:32]) - 1:0] EPCM;
	wire [$signed(P[4216-:32]) - 1:0] TrapVectorM;
	wire [1:0] MemRWE;
	wire [1:0] MemRWM;
	wire InstrValidD;
	wire InstrValidE;
	wire InstrValidM;
	wire InstrMisalignedFaultM;
	wire IllegalBaseInstrD;
	wire IllegalFPUInstrD;
	wire IllegalIEUFPUInstrD;
	wire InstrPageFaultF;
	wire LoadPageFaultM;
	wire StoreAmoPageFaultM;
	wire LoadMisalignedFaultM;
	wire LoadAccessFaultM;
	wire StoreAmoMisalignedFaultM;
	wire StoreAmoAccessFaultM;
	wire InvalidateICacheM;
	wire FlushDCacheM;
	wire PCSrcE;
	wire CSRWriteFenceM;
	wire DivBusyE;
	wire StructuralStallD;
	wire LoadStallD;
	wire StoreStallD;
	wire SquashSCW;
	wire MDUActiveE;
	wire ENVCFG_ADUE;
	wire ENVCFG_PBMTE;
	wire [3:0] ENVCFG_CBE;
	wire [3:0] CMOpM;
	wire IFUPrefetchE;
	wire LSUPrefetchM;
	wire [2:0] FRM_REGW;
	wire [4:0] RdE;
	wire [4:0] RdM;
	wire [4:0] RdW;
	wire FPUStallD;
	wire FWriteIntE;
	wire [$signed(P[901-:32]) - 1:0] FWriteDataM;
	wire [$signed(P[4216-:32]) - 1:0] FIntResM;
	wire [$signed(P[4216-:32]) - 1:0] FCvtIntResW;
	wire FCvtIntW;
	wire FDivBusyE;
	wire FRegWriteM;
	wire FpLoadStoreM;
	wire [4:0] SetFflagsM;
	wire [$signed(P[4216-:32]) - 1:0] FIntDivResultW;
	wire ITLBWriteF;
	wire ITLBMissOrUpdateAF;
	wire [$signed(P[4216-:32]) - 1:0] SATP_REGW;
	wire STATUS_MXR;
	wire STATUS_SUM;
	wire STATUS_MPRV;
	wire [1:0] STATUS_MPP;
	wire [1:0] STATUS_FS;
	wire [1:0] PrivilegeModeW;
	wire [$signed(P[4216-:32]) - 1:0] PTE;
	wire [1:0] PageType;
	wire sfencevmaM;
	wire SelHPTW;
	wire [(($signed(P[1640-:32]) - 3) >= 0 ? ($signed(P[3728-:32]) * ($signed(P[1640-:32]) - 2)) - 1 : ($signed(P[3728-:32]) * (4 - $signed(P[1640-:32]))) + ($signed(P[1640-:32]) - 4)):(($signed(P[1640-:32]) - 3) >= 0 ? 0 : $signed(P[1640-:32]) - 3)] PMPADDR_ARRAY_REGW;
	wire [($signed(P[3728-:32]) * 8) - 1:0] PMPCFG_ARRAY_REGW;
	wire IFUStallF;
	wire LSUStallM;
	wire [2:0] Funct3M;
	wire [$signed(P[4216-:32]) - 1:0] IEUAdrE;
	wire [$signed(P[4216-:32]) - 1:0] WriteDataM;
	wire [$signed(P[4216-:32]) - 1:0] IEUAdrM;
	wire [$signed(P[4216-:32]) - 1:0] IEUAdrxTvalM;
	wire [$signed(P[383-:32]) - 1:0] ReadDataW;
	wire CommittedM;
	wire [$signed(P[1640-:32]) - 1:0] IFUHADDR;
	wire [2:0] IFUHBURST;
	wire [1:0] IFUHTRANS;
	wire [2:0] IFUHSIZE;
	wire IFUHWRITE;
	wire IFUHREADY;
	wire [$signed(P[1640-:32]) - 1:0] LSUHADDR;
	wire [$signed(P[4216-:32]) - 1:0] LSUHWDATA;
	wire [($signed(P[4216-:32]) / 8) - 1:0] LSUHWSTRB;
	wire LSUHWRITE;
	wire LSUHREADY;
	wire BPWrongE;
	wire BPWrongM;
	wire BPDirWrongM;
	wire BTAWrongM;
	wire RASPredPCWrongM;
	wire IClassWrongM;
	wire [3:0] IClassM;
	wire InstrAccessFaultF;
	wire HPTWInstrAccessFaultF;
	wire HPTWInstrPageFaultF;
	wire [2:0] LSUHSIZE;
	wire [2:0] LSUHBURST;
	wire [1:0] LSUHTRANS;
	wire DCacheMiss;
	wire DCacheAccess;
	wire ICacheMiss;
	wire ICacheAccess;
	wire BigEndianM;
	wire FCvtIntE;
	wire CommittedF;
	wire BranchD;
	wire BranchE;
	wire JumpD;
	wire JumpE;
	wire DCacheStallM;
	wire ICacheStallF;
	wire wfiM;
	wire IntPendingM;
	ifu #(.P(P)) ifu(
		.clk(clk),
		.reset(reset),
		.StallF(StallF),
		.StallD(StallD),
		.StallE(StallE),
		.StallM(StallM),
		.StallW(StallW),
		.FlushD(FlushD),
		.FlushE(FlushE),
		.FlushM(FlushM),
		.FlushW(FlushW),
		.InstrValidE(InstrValidE),
		.InstrValidD(InstrValidD),
		.BranchD(BranchD),
		.BranchE(BranchE),
		.JumpD(JumpD),
		.JumpE(JumpE),
		.ICacheStallF(ICacheStallF),
		.HRDATA(HRDATA),
		.PCSpillF(PCSpillF),
		.IFUHADDR(IFUHADDR),
		.IFUStallF(IFUStallF),
		.IFUHBURST(IFUHBURST),
		.IFUHTRANS(IFUHTRANS),
		.IFUHSIZE(IFUHSIZE),
		.IFUHREADY(IFUHREADY),
		.IFUHWRITE(IFUHWRITE),
		.ICacheAccess(ICacheAccess),
		.ICacheMiss(ICacheMiss),
		.PCLinkE(PCLinkE),
		.PCSrcE(PCSrcE),
		.IEUAdrE(IEUAdrE),
		.IEUAdrM(IEUAdrM),
		.PCE(PCE),
		.BPWrongE(BPWrongE),
		.BPWrongM(BPWrongM),
		.CommittedF(CommittedF),
		.EPCM(EPCM),
		.TrapVectorM(TrapVectorM),
		.RetM(RetM),
		.TrapM(TrapM),
		.InvalidateICacheM(InvalidateICacheM),
		.CSRWriteFenceM(CSRWriteFenceM),
		.InstrD(InstrD),
		.InstrM(InstrM),
		.InstrOrigM(InstrOrigM),
		.PCM(PCM),
		.IClassM(IClassM),
		.BPDirWrongM(BPDirWrongM),
		.BTAWrongM(BTAWrongM),
		.RASPredPCWrongM(RASPredPCWrongM),
		.IClassWrongM(IClassWrongM),
		.IllegalBaseInstrD(IllegalBaseInstrD),
		.IllegalFPUInstrD(IllegalFPUInstrD),
		.InstrPageFaultF(InstrPageFaultF),
		.IllegalIEUFPUInstrD(IllegalIEUFPUInstrD),
		.InstrMisalignedFaultM(InstrMisalignedFaultM),
		.PrivilegeModeW(PrivilegeModeW),
		.PTE(PTE),
		.PageType(PageType),
		.SATP_REGW(SATP_REGW),
		.STATUS_MXR(STATUS_MXR),
		.STATUS_SUM(STATUS_SUM),
		.STATUS_MPRV(STATUS_MPRV),
		.STATUS_MPP(STATUS_MPP),
		.ENVCFG_PBMTE(ENVCFG_PBMTE),
		.ENVCFG_ADUE(ENVCFG_ADUE),
		.ITLBWriteF(ITLBWriteF),
		.sfencevmaM(sfencevmaM),
		.ITLBMissOrUpdateAF(ITLBMissOrUpdateAF),
		.PMPCFG_ARRAY_REGW(PMPCFG_ARRAY_REGW),
		.PMPADDR_ARRAY_REGW(PMPADDR_ARRAY_REGW),
		.InstrAccessFaultF(InstrAccessFaultF)
	);
	ieu #(.P(P)) ieu(
		.clk(clk),
		.reset(reset),
		.InstrD(InstrD),
		.STATUS_FS(STATUS_FS),
		.ENVCFG_CBE(ENVCFG_CBE),
		.IllegalIEUFPUInstrD(IllegalIEUFPUInstrD),
		.IllegalBaseInstrD(IllegalBaseInstrD),
		.PCE(PCE),
		.PCLinkE(PCLinkE),
		.FWriteIntE(FWriteIntE),
		.FCvtIntE(FCvtIntE),
		.IEUAdrE(IEUAdrE),
		.IntDivE(IntDivE),
		.W64E(W64E),
		.Funct3E(Funct3E),
		.ForwardedSrcAE(ForwardedSrcAE),
		.ForwardedSrcBE(ForwardedSrcBE),
		.MDUActiveE(MDUActiveE),
		.CMOpM(CMOpM),
		.IFUPrefetchE(IFUPrefetchE),
		.LSUPrefetchM(LSUPrefetchM),
		.SquashSCW(SquashSCW),
		.MemRWE(MemRWE),
		.MemRWM(MemRWM),
		.AtomicM(AtomicM),
		.WriteDataM(WriteDataM),
		.Funct3M(Funct3M),
		.SrcAM(SrcAM),
		.RdE(RdE),
		.RdM(RdM),
		.FIntResM(FIntResM),
		.FlushDCacheM(FlushDCacheM),
		.BranchD(BranchD),
		.BranchE(BranchE),
		.JumpD(JumpD),
		.JumpE(JumpE),
		.CSRReadValW(CSRReadValW),
		.MDUResultW(MDUResultW),
		.FIntDivResultW(FIntDivResultW),
		.RdW(RdW),
		.ReadDataW(ReadDataW[$signed(P[4216-:32]) - 1:0]),
		.InstrValidM(InstrValidM),
		.InstrValidE(InstrValidE),
		.InstrValidD(InstrValidD),
		.FCvtIntResW(FCvtIntResW),
		.FCvtIntW(FCvtIntW),
		.StallD(StallD),
		.StallE(StallE),
		.StallM(StallM),
		.StallW(StallW),
		.FlushD(FlushD),
		.FlushE(FlushE),
		.FlushM(FlushM),
		.FlushW(FlushW),
		.StructuralStallD(StructuralStallD),
		.LoadStallD(LoadStallD),
		.StoreStallD(StoreStallD),
		.PCSrcE(PCSrcE),
		.CSRReadM(CSRReadM),
		.CSRWriteM(CSRWriteM),
		.PrivilegedM(PrivilegedM),
		.CSRWriteFenceM(CSRWriteFenceM),
		.InvalidateICacheM(InvalidateICacheM)
	);
	lsu #(.P(P)) lsu(
		.clk(clk),
		.reset(reset),
		.StallM(StallM),
		.FlushM(FlushM),
		.StallW(StallW),
		.FlushW(FlushW),
		.MemRWE(MemRWE),
		.MemRWM(MemRWM),
		.Funct3M(Funct3M),
		.Funct7M(InstrM[31:25]),
		.AtomicM(AtomicM),
		.CommittedM(CommittedM),
		.DCacheMiss(DCacheMiss),
		.DCacheAccess(DCacheAccess),
		.SquashSCW(SquashSCW),
		.FpLoadStoreM(FpLoadStoreM),
		.FWriteDataM(FWriteDataM),
		.IEUAdrE(IEUAdrE),
		.IEUAdrM(IEUAdrM),
		.WriteDataM(WriteDataM),
		.ReadDataW(ReadDataW),
		.FlushDCacheM(FlushDCacheM),
		.CMOpM(CMOpM),
		.LSUPrefetchM(LSUPrefetchM),
		.LSUHADDR(LSUHADDR),
		.HRDATA(HRDATA),
		.LSUHWDATA(LSUHWDATA),
		.LSUHWSTRB(LSUHWSTRB),
		.LSUHSIZE(LSUHSIZE),
		.LSUHBURST(LSUHBURST),
		.LSUHTRANS(LSUHTRANS),
		.LSUHWRITE(LSUHWRITE),
		.LSUHREADY(LSUHREADY),
		.PrivilegeModeW(PrivilegeModeW),
		.BigEndianM(BigEndianM),
		.PMPCFG_ARRAY_REGW(PMPCFG_ARRAY_REGW),
		.PMPADDR_ARRAY_REGW(PMPADDR_ARRAY_REGW),
		.SATP_REGW(SATP_REGW),
		.STATUS_MXR(STATUS_MXR),
		.STATUS_SUM(STATUS_SUM),
		.STATUS_MPRV(STATUS_MPRV),
		.STATUS_MPP(STATUS_MPP),
		.ENVCFG_PBMTE(ENVCFG_PBMTE),
		.ENVCFG_ADUE(ENVCFG_ADUE),
		.sfencevmaM(sfencevmaM),
		.DCacheStallM(DCacheStallM),
		.IEUAdrxTvalM(IEUAdrxTvalM),
		.LoadPageFaultM(LoadPageFaultM),
		.StoreAmoPageFaultM(StoreAmoPageFaultM),
		.LoadMisalignedFaultM(LoadMisalignedFaultM),
		.LoadAccessFaultM(LoadAccessFaultM),
		.HPTWInstrAccessFaultF(HPTWInstrAccessFaultF),
		.HPTWInstrPageFaultF(HPTWInstrPageFaultF),
		.StoreAmoMisalignedFaultM(StoreAmoMisalignedFaultM),
		.StoreAmoAccessFaultM(StoreAmoAccessFaultM),
		.PCSpillF(PCSpillF),
		.ITLBMissOrUpdateAF(ITLBMissOrUpdateAF),
		.PTE(PTE),
		.PageType(PageType),
		.ITLBWriteF(ITLBWriteF),
		.SelHPTW(SelHPTW),
		.LSUStallM(LSUStallM)
	);
	generate
		if (P[4052]) begin : ebu
			ebu #(.P(P)) ebu(
				.clk(clk),
				.reset(reset),
				.IFUHADDR(IFUHADDR),
				.IFUHBURST(IFUHBURST),
				.IFUHTRANS(IFUHTRANS),
				.IFUHREADY(IFUHREADY),
				.IFUHSIZE(IFUHSIZE),
				.LSUHADDR(LSUHADDR),
				.LSUHWDATA(LSUHWDATA),
				.LSUHWSTRB(LSUHWSTRB),
				.LSUHSIZE(LSUHSIZE),
				.LSUHBURST(LSUHBURST),
				.LSUHTRANS(LSUHTRANS),
				.LSUHWRITE(LSUHWRITE),
				.LSUHREADY(LSUHREADY),
				.HREADY(HREADY),
				.HRESP(HRESP),
				.HCLK(HCLK),
				.HRESETn(HRESETn),
				.HADDR(HADDR),
				.HWDATA(HWDATA),
				.HWSTRB(HWSTRB),
				.HWRITE(HWRITE),
				.HSIZE(HSIZE),
				.HBURST(HBURST),
				.HPROT(HPROT),
				.HTRANS(HTRANS),
				.HMASTLOCK(HMASTLOCK)
			);
		end
		else begin : genblk1
			assign {IFUHREADY, LSUHREADY, HCLK, HRESETn, HADDR, HWDATA, HWSTRB, HWRITE, HSIZE, HBURST, HPROT, HTRANS, HMASTLOCK} = 1'sb0;
		end
	endgenerate
	hazard hzu(
		.BPWrongE(BPWrongE),
		.CSRWriteFenceM(CSRWriteFenceM),
		.RetM(RetM),
		.TrapM(TrapM),
		.StructuralStallD(StructuralStallD),
		.LSUStallM(LSUStallM),
		.IFUStallF(IFUStallF),
		.FPUStallD(FPUStallD),
		.ExternalStall(ExternalStall),
		.DivBusyE(DivBusyE),
		.FDivBusyE(FDivBusyE),
		.wfiM(wfiM),
		.IntPendingM(IntPendingM),
		.StallF(StallF),
		.StallD(StallD),
		.StallE(StallE),
		.StallM(StallM),
		.StallW(StallW),
		.FlushD(FlushD),
		.FlushE(FlushE),
		.FlushM(FlushM),
		.FlushW(FlushW)
	);
	generate
		if (P[4086]) begin : priv
			privileged #(.P(P)) priv(
				.clk(clk),
				.reset(reset),
				.FlushD(FlushD),
				.FlushE(FlushE),
				.FlushM(FlushM),
				.FlushW(FlushW),
				.StallD(StallD),
				.StallE(StallE),
				.StallM(StallM),
				.StallW(StallW),
				.CSRReadM(CSRReadM),
				.CSRWriteM(CSRWriteM),
				.SrcAM(SrcAM),
				.PCM(PCM),
				.InstrM(InstrM),
				.InstrOrigM(InstrOrigM),
				.CSRReadValW(CSRReadValW),
				.EPCM(EPCM),
				.TrapVectorM(TrapVectorM),
				.RetM(RetM),
				.TrapM(TrapM),
				.sfencevmaM(sfencevmaM),
				.InvalidateICacheM(InvalidateICacheM),
				.DCacheStallM(DCacheStallM),
				.ICacheStallF(ICacheStallF),
				.InstrValidM(InstrValidM),
				.CommittedM(CommittedM),
				.CommittedF(CommittedF),
				.FRegWriteM(FRegWriteM),
				.LoadStallD(LoadStallD),
				.StoreStallD(StoreStallD),
				.BPDirWrongM(BPDirWrongM),
				.BTAWrongM(BTAWrongM),
				.BPWrongM(BPWrongM),
				.RASPredPCWrongM(RASPredPCWrongM),
				.IClassWrongM(IClassWrongM),
				.DivBusyE(DivBusyE),
				.FDivBusyE(FDivBusyE),
				.IClassM(IClassM),
				.DCacheMiss(DCacheMiss),
				.DCacheAccess(DCacheAccess),
				.ICacheMiss(ICacheMiss),
				.ICacheAccess(ICacheAccess),
				.PrivilegedM(PrivilegedM),
				.InstrPageFaultF(InstrPageFaultF),
				.LoadPageFaultM(LoadPageFaultM),
				.StoreAmoPageFaultM(StoreAmoPageFaultM),
				.InstrMisalignedFaultM(InstrMisalignedFaultM),
				.IllegalIEUFPUInstrD(IllegalIEUFPUInstrD),
				.LoadMisalignedFaultM(LoadMisalignedFaultM),
				.StoreAmoMisalignedFaultM(StoreAmoMisalignedFaultM),
				.MTimerInt(MTimerInt),
				.MExtInt(MExtInt),
				.SExtInt(SExtInt),
				.MSwInt(MSwInt),
				.MTIME_CLINT(MTIME_CLINT),
				.IEUAdrxTvalM(IEUAdrxTvalM),
				.SetFflagsM(SetFflagsM),
				.InstrAccessFaultF(InstrAccessFaultF),
				.HPTWInstrAccessFaultF(HPTWInstrAccessFaultF),
				.HPTWInstrPageFaultF(HPTWInstrPageFaultF),
				.LoadAccessFaultM(LoadAccessFaultM),
				.StoreAmoAccessFaultM(StoreAmoAccessFaultM),
				.SelHPTW(SelHPTW),
				.PrivilegeModeW(PrivilegeModeW),
				.SATP_REGW(SATP_REGW),
				.STATUS_MXR(STATUS_MXR),
				.STATUS_SUM(STATUS_SUM),
				.STATUS_MPRV(STATUS_MPRV),
				.STATUS_MPP(STATUS_MPP),
				.STATUS_FS(STATUS_FS),
				.PMPCFG_ARRAY_REGW(PMPCFG_ARRAY_REGW),
				.PMPADDR_ARRAY_REGW(PMPADDR_ARRAY_REGW),
				.FRM_REGW(FRM_REGW),
				.ENVCFG_CBE(ENVCFG_CBE),
				.ENVCFG_PBMTE(ENVCFG_PBMTE),
				.ENVCFG_ADUE(ENVCFG_ADUE),
				.wfiM(wfiM),
				.IntPendingM(IntPendingM),
				.BigEndianM(BigEndianM)
			);
		end
		else begin : genblk2
			assign {CSRReadValW, PrivilegeModeW, SATP_REGW, STATUS_MXR, STATUS_SUM, STATUS_MPRV, STATUS_MPP, STATUS_FS, FRM_REGW, ENVCFG_CBE, ENVCFG_PBMTE, ENVCFG_ADUE, EPCM, TrapVectorM, RetM, TrapM, sfencevmaM, BigEndianM, wfiM, IntPendingM} = 1'sb0;
		end
		if (P[4063]) begin : mdu
			mdu #(.P(P)) mdu(
				.clk(clk),
				.reset(reset),
				.StallM(StallM),
				.StallW(StallW),
				.FlushE(FlushE),
				.FlushM(FlushM),
				.FlushW(FlushW),
				.ForwardedSrcAE(ForwardedSrcAE),
				.ForwardedSrcBE(ForwardedSrcBE),
				.Funct3E(Funct3E),
				.Funct3M(Funct3M),
				.IntDivE(IntDivE),
				.W64E(W64E),
				.MDUActiveE(MDUActiveE),
				.MDUResultW(MDUResultW),
				.DivBusyE(DivBusyE)
			);
		end
		else begin : genblk3
			assign MDUResultW = 1'sb0;
			assign DivBusyE = 1'b0;
		end
		if (P[1491]) begin : fpu
			fpu #(.P(P)) fpu(
				.clk(clk),
				.reset(reset),
				.FRM_REGW(FRM_REGW),
				.InstrD(InstrD),
				.ReadDataW(ReadDataW[$signed(P[901-:32]) - 1:0]),
				.ForwardedSrcAE(ForwardedSrcAE),
				.StallE(StallE),
				.StallM(StallM),
				.StallW(StallW),
				.FlushE(FlushE),
				.FlushM(FlushM),
				.FlushW(FlushW),
				.RdE(RdE),
				.RdM(RdM),
				.RdW(RdW),
				.STATUS_FS(STATUS_FS),
				.FRegWriteM(FRegWriteM),
				.FpLoadStoreM(FpLoadStoreM),
				.ForwardedSrcBE(ForwardedSrcBE),
				.Funct3E(Funct3E),
				.Funct3M(Funct3M),
				.IntDivE(IntDivE),
				.W64E(W64E),
				.FPUStallD(FPUStallD),
				.FWriteIntE(FWriteIntE),
				.FCvtIntE(FCvtIntE),
				.FWriteDataM(FWriteDataM),
				.FIntResM(FIntResM),
				.FCvtIntResW(FCvtIntResW),
				.FCvtIntW(FCvtIntW),
				.FDivBusyE(FDivBusyE),
				.IllegalFPUInstrD(IllegalFPUInstrD),
				.SetFflagsM(SetFflagsM),
				.FIntDivResultW(FIntDivResultW)
			);
		end
		else begin : genblk4
			assign {FPUStallD, FWriteIntE, FCvtIntE, FIntResM, FCvtIntW, FRegWriteM, IllegalFPUInstrD, SetFflagsM, FpLoadStoreM, FWriteDataM, FCvtIntResW, FIntDivResultW, FDivBusyE} = 1'sb0;
		end
	endgenerate
endmodule
module wallypipelinedsoc (
	clk,
	reset_ext,
	reset,
	HRDATAEXT,
	HREADYEXT,
	HRESPEXT,
	HSELEXT,
	ExternalStall,
	HCLK,
	HRESETn,
	HADDR,
	HWDATA,
	HWSTRB,
	HWRITE,
	HSIZE,
	HBURST,
	HPROT,
	HTRANS,
	HMASTLOCK,
	HREADY,
	TIMECLK,
	GPIOIN,
	GPIOOUT,
	GPIOEN,
	UARTSin,
	UARTSout,
	SPIIn,
	SPIOut,
	SPICS,
	SPICLK,
	SDCIn,
	SDCCmd,
	SDCCS,
	SDCCLK
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset_ext;
	output wire reset;
	input wire [$signed(P[4151-:32]) - 1:0] HRDATAEXT;
	input wire HREADYEXT;
	input wire HRESPEXT;
	output wire HSELEXT;
	input wire ExternalStall;
	output wire HCLK;
	output wire HRESETn;
	output wire [$signed(P[1640-:32]) - 1:0] HADDR;
	output wire [$signed(P[4151-:32]) - 1:0] HWDATA;
	output wire [($signed(P[4216-:32]) / 8) - 1:0] HWSTRB;
	output wire HWRITE;
	output wire [2:0] HSIZE;
	output wire [2:0] HBURST;
	output wire [3:0] HPROT;
	output wire [1:0] HTRANS;
	output wire HMASTLOCK;
	output wire HREADY;
	input wire TIMECLK;
	input wire [31:0] GPIOIN;
	output wire [31:0] GPIOOUT;
	output wire [31:0] GPIOEN;
	input wire UARTSin;
	output wire UARTSout;
	input wire SPIIn;
	output wire SPIOut;
	output wire [3:0] SPICS;
	output wire SPICLK;
	input wire SDCIn;
	output wire SDCCmd;
	output wire [3:0] SDCCS;
	output wire SDCCLK;
	wire [$signed(P[4151-:32]) - 1:0] HRDATA;
	wire HRESP;
	wire MTimerInt;
	wire MSwInt;
	wire [63:0] MTIME_CLINT;
	wire MExtInt;
	wire SExtInt;
	synchronizer resetsync(
		.clk(clk),
		.d(reset_ext),
		.q(reset)
	);
	wallypipelinedcore #(.P(P)) core(
		.clk(clk),
		.reset(reset),
		.MTimerInt(MTimerInt),
		.MExtInt(MExtInt),
		.SExtInt(SExtInt),
		.MSwInt(MSwInt),
		.MTIME_CLINT(MTIME_CLINT),
		.HRDATA(HRDATA),
		.HREADY(HREADY),
		.HRESP(HRESP),
		.HCLK(HCLK),
		.HRESETn(HRESETn),
		.HADDR(HADDR),
		.HWDATA(HWDATA),
		.HWSTRB(HWSTRB),
		.HWRITE(HWRITE),
		.HSIZE(HSIZE),
		.HBURST(HBURST),
		.HPROT(HPROT),
		.HTRANS(HTRANS),
		.HMASTLOCK(HMASTLOCK),
		.ExternalStall(ExternalStall)
	);
	generate
		if (P[4052]) begin : uncoregen
			uncore #(.P(P)) uncore(
				.HCLK(HCLK),
				.HRESETn(HRESETn),
				.TIMECLK(TIMECLK),
				.HADDR(HADDR),
				.HWDATA(HWDATA),
				.HWSTRB(HWSTRB),
				.HWRITE(HWRITE),
				.HSIZE(HSIZE),
				.HBURST(HBURST),
				.HPROT(HPROT),
				.HTRANS(HTRANS),
				.HMASTLOCK(HMASTLOCK),
				.HRDATAEXT(HRDATAEXT),
				.HREADYEXT(HREADYEXT),
				.HRESPEXT(HRESPEXT),
				.HRDATA(HRDATA),
				.HREADY(HREADY),
				.HRESP(HRESP),
				.HSELEXT(HSELEXT),
				.MTimerInt(MTimerInt),
				.MSwInt(MSwInt),
				.MExtInt(MExtInt),
				.SExtInt(SExtInt),
				.GPIOIN(GPIOIN),
				.GPIOOUT(GPIOOUT),
				.GPIOEN(GPIOEN),
				.UARTSin(UARTSin),
				.UARTSout(UARTSout),
				.MTIME_CLINT(MTIME_CLINT),
				.SPIIn(SPIIn),
				.SPIOut(SPIOut),
				.SPICS(SPICS),
				.SPICLK(SPICLK),
				.SDCIn(SDCIn),
				.SDCCmd(SDCCmd),
				.SDCCS(SDCCS),
				.SDCCLK(SDCCLK)
			);
		end
		else begin : genblk1
			assign {HRDATA, HREADY, HRESP, HSELEXT, MTimerInt, MSwInt, MExtInt, SExtInt, MTIME_CLINT, GPIOOUT, GPIOEN, UARTSout, SPIOut, SPICS, SPICLK, SDCCmd, SDCCS, SDCCLK} = 1'sb0;
		end
	endgenerate
endmodule
module fdivsqrt (
	clk,
	reset,
	FmtE,
	XsE,
	XmE,
	YmE,
	XeE,
	YeE,
	XInfE,
	YInfE,
	XZeroE,
	YZeroE,
	XNaNE,
	YNaNE,
	BiasE,
	NfE,
	FDivStartE,
	IDivStartE,
	StallM,
	FlushE,
	SqrtE,
	SqrtM,
	ForwardedSrcAE,
	ForwardedSrcBE,
	Funct3E,
	Funct3M,
	IntDivE,
	W64E,
	DivStickyM,
	FDivBusyE,
	IFDivStartE,
	FDivDoneE,
	UeM,
	UmM,
	FIntDivResultM
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire [$signed(P[707-:32]) - 1:0] FmtE;
	input wire XsE;
	input wire [$signed(P[805-:32]):0] XmE;
	input wire [$signed(P[805-:32]):0] YmE;
	input wire [$signed(P[837-:32]) - 1:0] XeE;
	input wire [$signed(P[837-:32]) - 1:0] YeE;
	input wire XInfE;
	input wire YInfE;
	input wire XZeroE;
	input wire YZeroE;
	input wire XNaNE;
	input wire YNaNE;
	input wire [$signed(P[837-:32]) - 2:0] BiasE;
	input wire [$signed(P[869-:32]) - 1:0] NfE;
	input wire FDivStartE;
	input wire IDivStartE;
	input wire StallM;
	input wire FlushE;
	input wire SqrtE;
	input wire SqrtM;
	input wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcAE;
	input wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcBE;
	input wire [2:0] Funct3E;
	input wire [2:0] Funct3M;
	input wire IntDivE;
	input wire W64E;
	output wire DivStickyM;
	output wire FDivBusyE;
	output wire IFDivStartE;
	output wire FDivDoneE;
	output wire [$signed(P[837-:32]) + 1:0] UeM;
	output wire [$signed(P[95-:32]):0] UmM;
	output wire [$signed(P[4216-:32]) - 1:0] FIntDivResultM;
	wire [$signed(P[95-:32]) + 3:0] WS;
	wire [$signed(P[95-:32]) + 3:0] WC;
	wire [$signed(P[95-:32]) + 3:0] X;
	wire [$signed(P[95-:32]) + 3:0] D;
	wire [$signed(P[95-:32]):0] FirstU;
	wire [$signed(P[95-:32]):0] FirstUM;
	wire [$signed(P[95-:32]) + 1:0] FirstC;
	wire WZeroE;
	wire [$signed(P[127-:32]) - 1:0] CyclesE;
	wire SpecialCaseM;
	wire BZeroM;
	wire [$signed(P[63-:32]) - 1:0] IntNormShiftM;
	wire ALTBM;
	wire AsM;
	wire BsM;
	wire W64M;
	wire [$signed(P[4216-:32]) - 1:0] AM;
	wire ISpecialCaseE;
	fdivsqrtpreproc #(.P(P)) fdivsqrtpreproc(
		.clk(clk),
		.IFDivStartE(IFDivStartE),
		.Xm(XmE),
		.Ym(YmE),
		.Xe(XeE),
		.Ye(YeE),
		.FmtE(FmtE),
		.Bias(BiasE),
		.Nf(NfE),
		.SqrtE(SqrtE),
		.XZeroE(XZeroE),
		.Funct3E(Funct3E),
		.UeM(UeM),
		.X(X),
		.D(D),
		.CyclesE(CyclesE),
		.ForwardedSrcAE(ForwardedSrcAE),
		.ForwardedSrcBE(ForwardedSrcBE),
		.IntDivE(IntDivE),
		.W64E(W64E),
		.ISpecialCaseE(ISpecialCaseE),
		.BZeroM(BZeroM),
		.IntNormShiftM(IntNormShiftM),
		.AM(AM),
		.W64M(W64M),
		.ALTBM(ALTBM),
		.AsM(AsM),
		.BsM(BsM)
	);
	fdivsqrtfsm #(.P(P)) fdivsqrtfsm(
		.clk(clk),
		.reset(reset),
		.XInfE(XInfE),
		.YInfE(YInfE),
		.XZeroE(XZeroE),
		.YZeroE(YZeroE),
		.XNaNE(XNaNE),
		.YNaNE(YNaNE),
		.FDivStartE(FDivStartE),
		.XsE(XsE),
		.SqrtE(SqrtE),
		.WZeroE(WZeroE),
		.FlushE(FlushE),
		.StallM(StallM),
		.FDivBusyE(FDivBusyE),
		.IFDivStartE(IFDivStartE),
		.FDivDoneE(FDivDoneE),
		.SpecialCaseM(SpecialCaseM),
		.CyclesE(CyclesE),
		.IDivStartE(IDivStartE),
		.ISpecialCaseE(ISpecialCaseE),
		.IntDivE(IntDivE)
	);
	fdivsqrtiter #(.P(P)) fdivsqrtiter(
		.clk(clk),
		.IFDivStartE(IFDivStartE),
		.FDivBusyE(FDivBusyE),
		.SqrtE(SqrtE),
		.X(X),
		.D(D),
		.FirstU(FirstU),
		.FirstUM(FirstUM),
		.FirstC(FirstC),
		.FirstWS(WS),
		.FirstWC(WC)
	);
	fdivsqrtpostproc #(.P(P)) fdivsqrtpostproc(
		.clk(clk),
		.reset(reset),
		.StallM(StallM),
		.WS(WS),
		.WC(WC),
		.D(D),
		.FirstU(FirstU),
		.FirstUM(FirstUM),
		.FirstC(FirstC),
		.SqrtE(SqrtE),
		.SqrtM(SqrtM),
		.SpecialCaseM(SpecialCaseM),
		.UmM(UmM),
		.WZeroE(WZeroE),
		.DivStickyM(DivStickyM),
		.IntNormShiftM(IntNormShiftM),
		.ALTBM(ALTBM),
		.AsM(AsM),
		.BsM(BsM),
		.BZeroM(BZeroM),
		.W64M(W64M),
		.RemOpM(Funct3M[1]),
		.AM(AM),
		.FIntDivResultM(FIntDivResultM)
	);
endmodule
module fdivsqrtcycles (
	Nf,
	IntDivE,
	IntResultBitsE,
	CyclesE
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[869-:32]) - 1:0] Nf;
	input wire IntDivE;
	input wire [$signed(P[63-:32]) - 1:0] IntResultBitsE;
	output reg [$signed(P[127-:32]) - 1:0] CyclesE;
	reg [$signed(P[63-:32]) - 1:0] FPResultBitsE;
	reg [$signed(P[63-:32]) - 1:0] ResultBitsE;
	always @(*) begin
		if (_sv2v_0)
			;
		FPResultBitsE = (Nf + 2) + $signed(P[223-:32]);
		if (P[3729])
			ResultBitsE = (IntDivE ? IntResultBitsE : FPResultBitsE);
		else
			ResultBitsE = FPResultBitsE;
		CyclesE = ((ResultBitsE - 1) / $signed(P[191-:32])) + 1;
	end
	initial _sv2v_0 = 0;
endmodule
module fdivsqrtexpcalc (
	Bias,
	Xe,
	Ye,
	Sqrt,
	ell,
	m,
	Ue
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[837-:32]) - 2:0] Bias;
	input wire [$signed(P[837-:32]) - 1:0] Xe;
	input wire [$signed(P[837-:32]) - 1:0] Ye;
	input wire Sqrt;
	input wire [$signed(P[63-:32]) - 1:0] ell;
	input wire [$signed(P[63-:32]) - 1:0] m;
	output wire [$signed(P[837-:32]) + 1:0] Ue;
	wire [$signed(P[837-:32]) + 1:0] SXExp;
	wire [$signed(P[837-:32]) + 1:0] SExp;
	wire [$signed(P[837-:32]) + 1:0] DExp;
	function automatic signed [(($signed(P[837-:32]) + 1) >= 0 ? $signed(P[837-:32]) + 2 : 1 - ($signed(P[837-:32]) + 1)) - 1:0] sv2v_cast_A1EFF_signed;
		input reg signed [(($signed(P[837-:32]) + 1) >= 0 ? $signed(P[837-:32]) + 2 : 1 - ($signed(P[837-:32]) + 1)) - 1:0] inp;
		sv2v_cast_A1EFF_signed = inp;
	endfunction
	assign SXExp = ({2'b00, Xe} - {{($signed(P[837-:32]) + 1) - $signed(P[63-:32]) {1'b0}}, ell}) - sv2v_cast_A1EFF_signed($signed(P[771-:32]));
	assign SExp = {SXExp[$signed(P[837-:32]) + 1], SXExp[$signed(P[837-:32]) + 1:1]} + {2'b00, Bias};
	assign DExp = ((({2'b00, Xe} - {{($signed(P[837-:32]) + 1) - $signed(P[63-:32]) {1'b0}}, ell}) - {2'b00, Ye}) + {{($signed(P[837-:32]) + 1) - $signed(P[63-:32]) {1'b0}}, m}) + {3'b000, Bias};
	assign Ue = (Sqrt ? SExp : DExp);
endmodule
module fdivsqrtfgen2 (
	up,
	uz,
	C,
	U,
	UM,
	F
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire up;
	input wire uz;
	input wire [$signed(P[95-:32]) + 3:0] C;
	input wire [$signed(P[95-:32]) + 3:0] U;
	input wire [$signed(P[95-:32]) + 3:0] UM;
	output reg [$signed(P[95-:32]) + 3:0] F;
	wire [$signed(P[95-:32]) + 3:0] FP;
	wire [$signed(P[95-:32]) + 3:0] FN;
	wire [$signed(P[95-:32]) + 3:0] FZ;
	assign FP = ~(U << 1) & C;
	assign FN = (UM << 1) | (C & ~(C << 2));
	assign FZ = 1'sb0;
	always @(*) begin
		if (_sv2v_0)
			;
		if (up)
			F = FP;
		else if (uz)
			F = FZ;
		else
			F = FN;
	end
	initial _sv2v_0 = 0;
endmodule
module fdivsqrtfgen4 (
	udigit,
	C,
	U,
	UM,
	F
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [3:0] udigit;
	input wire [$signed(P[95-:32]) + 3:0] C;
	input wire [$signed(P[95-:32]) + 3:0] U;
	input wire [$signed(P[95-:32]) + 3:0] UM;
	output reg [$signed(P[95-:32]) + 3:0] F;
	wire [$signed(P[95-:32]) + 3:0] F2;
	wire [$signed(P[95-:32]) + 3:0] F1;
	wire [$signed(P[95-:32]) + 3:0] F0;
	wire [$signed(P[95-:32]) + 3:0] FN1;
	wire [$signed(P[95-:32]) + 3:0] FN2;
	assign F2 = (~U << 2) & (C << 2);
	assign F1 = ~(U << 1) & C;
	assign F0 = 1'sb0;
	assign FN1 = (UM << 1) | (C & ~(C << 3));
	assign FN2 = (UM << 2) | ((C << 2) & ~(C << 4));
	always @(*) begin
		if (_sv2v_0)
			;
		if (udigit[3])
			F = F2;
		else if (udigit[2])
			F = F1;
		else if (udigit[1])
			F = FN1;
		else if (udigit[0])
			F = FN2;
		else
			F = F0;
	end
	initial _sv2v_0 = 0;
endmodule
module fdivsqrtfsm (
	clk,
	reset,
	XInfE,
	YInfE,
	XZeroE,
	YZeroE,
	XNaNE,
	YNaNE,
	FDivStartE,
	IDivStartE,
	XsE,
	WZeroE,
	SqrtE,
	StallM,
	FlushE,
	IntDivE,
	ISpecialCaseE,
	CyclesE,
	IFDivStartE,
	FDivBusyE,
	FDivDoneE,
	SpecialCaseM
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire XInfE;
	input wire YInfE;
	input wire XZeroE;
	input wire YZeroE;
	input wire XNaNE;
	input wire YNaNE;
	input wire FDivStartE;
	input wire IDivStartE;
	input wire XsE;
	input wire WZeroE;
	input wire SqrtE;
	input wire StallM;
	input wire FlushE;
	input wire IntDivE;
	input wire ISpecialCaseE;
	input wire [$signed(P[127-:32]) - 1:0] CyclesE;
	output wire IFDivStartE;
	output wire FDivBusyE;
	output wire FDivDoneE;
	output wire SpecialCaseM;
	reg [1:0] state;
	wire SpecialCaseE;
	wire FSpecialCaseE;
	reg [$signed(P[127-:32]) - 1:0] step;
	assign IFDivStartE = ((FDivStartE | (IDivStartE & P[3729])) & (state == 2'd0)) & ~StallM;
	assign FDivDoneE = state == 2'd2;
	assign FDivBusyE = (state == 2'd1) | IFDivStartE;
	assign FSpecialCaseE = (((XZeroE | XInfE) | XNaNE) | (XsE & SqrtE)) | (((YZeroE | YInfE) | YNaNE) & ~SqrtE);
	generate
		if (P[3729]) begin : genblk1
			assign SpecialCaseE = (IntDivE ? ISpecialCaseE : FSpecialCaseE);
		end
		else begin : genblk1
			assign SpecialCaseE = FSpecialCaseE;
		end
	endgenerate
	flopenr #(.WIDTH(1)) SpecialCaseReg(
		.clk(clk),
		.reset(reset),
		.en(IFDivStartE),
		.d(SpecialCaseE),
		.q(SpecialCaseM)
	);
	always @(posedge clk)
		if (reset | FlushE)
			state <= 2'd0;
		else if (IFDivStartE) begin
			step <= CyclesE;
			if (SpecialCaseE)
				state <= 2'd2;
			else
				state <= 2'd1;
		end
		else if (state == 2'd1) begin
			if ((step == 1) | WZeroE)
				state <= 2'd2;
			step <= step - 1;
		end
		else if (state == 2'd2) begin
			if (StallM)
				state <= 2'd2;
			else
				state <= 2'd0;
		end
endmodule
module fdivsqrtiter (
	clk,
	IFDivStartE,
	FDivBusyE,
	SqrtE,
	X,
	D,
	FirstU,
	FirstUM,
	FirstC,
	FirstWS,
	FirstWC
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire IFDivStartE;
	input wire FDivBusyE;
	input wire SqrtE;
	input wire [$signed(P[95-:32]) + 3:0] X;
	input wire [$signed(P[95-:32]) + 3:0] D;
	output wire [$signed(P[95-:32]):0] FirstU;
	output wire [$signed(P[95-:32]):0] FirstUM;
	output wire [$signed(P[95-:32]) + 1:0] FirstC;
	output wire [$signed(P[95-:32]) + 3:0] FirstWS;
	output wire [$signed(P[95-:32]) + 3:0] FirstWC;
	wire [$signed(P[95-:32]) + 3:0] WSNext [$signed(P[1790-:32]) - 1:0];
	wire [$signed(P[95-:32]) + 3:0] WCNext [$signed(P[1790-:32]) - 1:0];
	wire [$signed(P[95-:32]) + 3:0] WS [$signed(P[1790-:32]):0];
	wire [$signed(P[95-:32]) + 3:0] WC [$signed(P[1790-:32]):0];
	wire [$signed(P[95-:32]):0] U [$signed(P[1790-:32]):0];
	wire [$signed(P[95-:32]):0] UM [$signed(P[1790-:32]):0];
	wire [$signed(P[95-:32]):0] UNext [$signed(P[1790-:32]) - 1:0];
	wire [$signed(P[95-:32]):0] UMNext [$signed(P[1790-:32]) - 1:0];
	wire [$signed(P[95-:32]) + 1:0] C [$signed(P[1790-:32]):0];
	wire [$signed(P[95-:32]) + 1:0] initC;
	wire [$signed(P[1790-:32]) - 1:0] un;
	wire [$signed(P[95-:32]) + 3:0] WSN;
	wire [$signed(P[95-:32]) + 3:0] WCN;
	wire [$signed(P[95-:32]) + 3:0] DBar;
	wire [$signed(P[95-:32]) + 3:0] D2;
	wire [$signed(P[95-:32]) + 3:0] DBar2;
	wire [$signed(P[95-:32]) + 1:0] NextC;
	wire [$signed(P[95-:32]):0] UMux;
	wire [$signed(P[95-:32]):0] UMMux;
	wire [$signed(P[95-:32]):0] initU;
	wire [$signed(P[95-:32]):0] initUM;
	mux2 #(.WIDTH($signed(P[95-:32]) + 4)) wsmux(
		.d0(WS[$signed(P[1790-:32])]),
		.d1(X),
		.s(IFDivStartE),
		.y(WSN)
	);
	localparam sv2v_uu_wcmux_WIDTH = $signed(P[95-:32]) + 4;
	localparam [sv2v_uu_wcmux_WIDTH - 1:0] sv2v_uu_wcmux_ext_d1_0 = 1'sb0;
	mux2 #(.WIDTH($signed(P[95-:32]) + 4)) wcmux(
		.d0(WC[$signed(P[1790-:32])]),
		.d1(sv2v_uu_wcmux_ext_d1_0),
		.s(IFDivStartE),
		.y(WCN)
	);
	flopen #(.WIDTH($signed(P[95-:32]) + 4)) wsreg(
		.clk(clk),
		.en(FDivBusyE),
		.d(WSN),
		.q(WS[0])
	);
	flopen #(.WIDTH($signed(P[95-:32]) + 4)) wcreg(
		.clk(clk),
		.en(FDivBusyE),
		.d(WCN),
		.q(WC[0])
	);
	assign initU = {$signed(P[95-:32]) + 1 {1'b0}};
	assign initUM = {1'b1, {$signed(P[95-:32]) {1'b0}}};
	mux2 #(.WIDTH($signed(P[95-:32]) + 1)) Umux(
		.d0(UNext[$signed(P[1790-:32]) - 1]),
		.d1(initU),
		.s(IFDivStartE),
		.y(UMux)
	);
	mux2 #(.WIDTH($signed(P[95-:32]) + 1)) UMmux(
		.d0(UMNext[$signed(P[1790-:32]) - 1]),
		.d1(initUM),
		.s(IFDivStartE),
		.y(UMMux)
	);
	flopen #(.WIDTH($signed(P[95-:32]) + 1)) UReg(
		.clk(clk),
		.en(FDivBusyE),
		.d(UMux),
		.q(U[0])
	);
	flopen #(.WIDTH($signed(P[95-:32]) + 1)) UMReg(
		.clk(clk),
		.en(FDivBusyE),
		.d(UMMux),
		.q(UM[0])
	);
	generate
		if ($signed(P[1822-:32]) == 4) begin : genblk1
			assign initC = 1'sb0;
		end
		else begin : genblk1
			assign initC = {2'b10, {$signed(P[95-:32]) {1'b0}}};
		end
	endgenerate
	mux2 #(.WIDTH($signed(P[95-:32]) + 2)) cmux(
		.d0(C[$signed(P[1790-:32])]),
		.d1(initC),
		.s(IFDivStartE),
		.y(NextC)
	);
	flopen #(.WIDTH($signed(P[95-:32]) + 2)) creg(
		.clk(clk),
		.en(FDivBusyE),
		.d(NextC),
		.q(C[0])
	);
	assign DBar = ~D;
	generate
		if ($signed(P[1822-:32]) == 4) begin : d2
			assign D2 = D << 1;
			assign DBar2 = ~D2;
		end
	endgenerate
	genvar _gv_i_7;
	generate
		for (_gv_i_7 = 0; $unsigned(_gv_i_7) < $signed(P[1790-:32]); _gv_i_7 = _gv_i_7 + 1) begin : iterations
			localparam i = _gv_i_7;
			if ($signed(P[1822-:32]) == 2) begin : stage
				fdivsqrtstage2 #(.P(P)) fdivsqrtstage(
					.D(D),
					.DBar(DBar),
					.SqrtE(SqrtE),
					.WS(WS[i]),
					.WC(WC[i]),
					.WSNext(WSNext[i]),
					.WCNext(WCNext[i]),
					.C(C[i]),
					.U(U[i]),
					.UM(UM[i]),
					.CNext(C[i + 1]),
					.UNext(UNext[i]),
					.UMNext(UMNext[i]),
					.un(un[i])
				);
			end
			else begin : stage
				fdivsqrtstage4 #(.P(P)) fdivsqrtstage(
					.D(D),
					.DBar(DBar),
					.D2(D2),
					.DBar2(DBar2),
					.SqrtE(SqrtE),
					.WS(WS[i]),
					.WC(WC[i]),
					.WSNext(WSNext[i]),
					.WCNext(WCNext[i]),
					.C(C[i]),
					.U(U[i]),
					.UM(UM[i]),
					.CNext(C[i + 1]),
					.UNext(UNext[i]),
					.UMNext(UMNext[i]),
					.un(un[i])
				);
			end
			assign WS[i + 1] = WSNext[i];
			assign WC[i + 1] = WCNext[i];
			assign U[i + 1] = UNext[i];
			assign UM[i + 1] = UMNext[i];
		end
	endgenerate
	assign FirstWS = WS[0];
	assign FirstWC = WC[0];
	assign FirstU = U[0];
	assign FirstUM = UM[0];
	assign FirstC = C[0];
endmodule
module fdivsqrtpostproc (
	clk,
	reset,
	StallM,
	WS,
	WC,
	D,
	FirstU,
	FirstUM,
	FirstC,
	SqrtE,
	SqrtM,
	SpecialCaseM,
	AM,
	RemOpM,
	ALTBM,
	BZeroM,
	AsM,
	BsM,
	W64M,
	IntNormShiftM,
	UmM,
	WZeroE,
	DivStickyM,
	FIntDivResultM
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallM;
	input wire [$signed(P[95-:32]) + 3:0] WS;
	input wire [$signed(P[95-:32]) + 3:0] WC;
	input wire [$signed(P[95-:32]) + 3:0] D;
	input wire [$signed(P[95-:32]):0] FirstU;
	input wire [$signed(P[95-:32]):0] FirstUM;
	input wire [$signed(P[95-:32]) + 1:0] FirstC;
	input wire SqrtE;
	input wire SqrtM;
	input wire SpecialCaseM;
	input wire [$signed(P[4216-:32]) - 1:0] AM;
	input wire RemOpM;
	input wire ALTBM;
	input wire BZeroM;
	input wire AsM;
	input wire BsM;
	input wire W64M;
	input wire [$signed(P[63-:32]) - 1:0] IntNormShiftM;
	output wire [$signed(P[95-:32]):0] UmM;
	output wire WZeroE;
	output wire DivStickyM;
	output wire [$signed(P[4216-:32]) - 1:0] FIntDivResultM;
	wire [$signed(P[95-:32]) + 3:0] Sum;
	wire [$signed(P[31-:32]) + 3:0] W;
	wire [$signed(P[95-:32]):0] PreUmM;
	wire NegStickyM;
	wire weq0E;
	wire WZeroM;
	reg [$signed(P[4216-:32]) - 1:0] IntDivResultM;
	wire NegQuotM;
	aplusbeq0 #(.WIDTH($signed(P[95-:32]) + 4)) wspluswceq0(
		.a(WS),
		.b(WC),
		.zero(weq0E)
	);
	generate
		if ($signed(P[1822-:32]) == 2) begin : R2EarlyTerm
			wire [$signed(P[95-:32]) + 3:0] FZeroE;
			wire [$signed(P[95-:32]) + 3:0] FZeroSqrtE;
			wire [$signed(P[95-:32]) + 3:0] FZeroDivE;
			wire [$signed(P[95-:32]) + 2:0] FirstK;
			wire wfeq0E;
			wire [$signed(P[95-:32]) + 3:0] WCF;
			wire [$signed(P[95-:32]) + 3:0] WSF;
			assign FirstK = {1'b1, FirstC} & ~({1'b1, FirstC} << 1);
			assign FZeroSqrtE = {FirstUM[$signed(P[95-:32])], FirstUM, 2'b00} | {FirstK, 1'b0};
			assign FZeroDivE = D << 1;
			mux2 #(.WIDTH($signed(P[95-:32]) + 4)) fzeromux(
				.d0(FZeroDivE),
				.d1(FZeroSqrtE),
				.s(SqrtE),
				.y(FZeroE)
			);
			csa #(.N($signed(P[95-:32]) + 4)) fadd(
				.x(WS),
				.y(WC),
				.z(FZeroE),
				.cin(1'b0),
				.s(WSF),
				.c(WCF)
			);
			aplusbeq0 #(.WIDTH($signed(P[95-:32]) + 4)) wcfpluswsfeq0(
				.a(WCF),
				.b(WSF),
				.zero(wfeq0E)
			);
			assign WZeroE = weq0E | wfeq0E;
		end
		else begin : genblk1
			assign WZeroE = weq0E;
		end
	endgenerate
	flopenr #(.WIDTH(1)) WZeroMReg(
		.clk(clk),
		.reset(reset),
		.en(~StallM),
		.d(WZeroE),
		.q(WZeroM)
	);
	assign DivStickyM = ~WZeroM & ~SpecialCaseM;
	assign Sum = WC + WS;
	assign NegStickyM = Sum[$signed(P[95-:32]) + 3];
	mux2 #(.WIDTH($signed(P[95-:32]) + 1)) preummux(
		.d0(FirstU),
		.d1(FirstUM),
		.s(NegStickyM),
		.y(PreUmM)
	);
	mux2 #(.WIDTH($signed(P[95-:32]) + 1)) ummux(
		.d0(PreUmM),
		.d1(PreUmM << 1),
		.s(SqrtM),
		.y(UmM)
	);
	generate
		if (P[3729]) begin : intpostproc
			wire [$signed(P[31-:32]) + 3:0] UnsignedQuotM;
			wire [$signed(P[31-:32]) + 3:0] NormRemM;
			wire [$signed(P[31-:32]) + 3:0] NormRemDM;
			wire [$signed(P[31-:32]) + 3:0] NormQuotM;
			wire signed [$signed(P[31-:32]) + 3:0] PreResultM;
			wire signed [$signed(P[31-:32]) + 3:0] PreResultShiftedM;
			wire signed [$signed(P[31-:32]) + 3:0] PreIntResultM;
			wire [$signed(P[31-:32]) + 3:0] DTrunc;
			wire [$signed(P[31-:32]) + 3:0] SumTrunc;
			assign SumTrunc = Sum[$signed(P[95-:32]) + 3:$signed(P[95-:32]) - $signed(P[31-:32])];
			assign DTrunc = D[$signed(P[95-:32]) + 3:$signed(P[95-:32]) - $signed(P[31-:32])];
			assign W = $signed(SumTrunc) >>> $signed(P[223-:32]);
			assign UnsignedQuotM = {3'b000, PreUmM[$signed(P[95-:32]):$signed(P[95-:32]) - $signed(P[31-:32])]};
			assign NegQuotM = AsM ^ BsM;
			mux2 #(.WIDTH($signed(P[31-:32]) + 4)) normremdmux(
				.d0(W),
				.d1(W + DTrunc),
				.s(NegStickyM),
				.y(NormRemDM)
			);
			mux2 #(.WIDTH($signed(P[31-:32]) + 4)) presresultmux(
				.d0(UnsignedQuotM),
				.d1(NormRemDM),
				.s(RemOpM),
				.y(PreResultM)
			);
			assign PreResultShiftedM = PreResultM >> IntNormShiftM;
			mux2 #(.WIDTH($signed(P[31-:32]) + 4)) preintresultmux(
				.d0(PreResultShiftedM),
				.d1(-PreResultShiftedM),
				.s(AsM ^ (BsM & ~RemOpM)),
				.y(PreIntResultM)
			);
			always @(*) begin
				if (_sv2v_0)
					;
				if (BZeroM) begin
					if (RemOpM)
						IntDivResultM = AM;
					else
						IntDivResultM = {$signed(P[4216-:32]) {1'b1}};
				end
				else if (ALTBM) begin
					if (RemOpM)
						IntDivResultM = AM;
					else
						IntDivResultM = 1'sb0;
				end
				else
					IntDivResultM = PreIntResultM[$signed(P[4216-:32]) - 1:0];
			end
			if ($signed(P[4216-:32]) == 64) begin : genblk1
				mux2 #(.WIDTH(64)) resmux(
					.d0(IntDivResultM[$signed(P[4216-:32]) - 1:0]),
					.d1({{$signed(P[4216-:32]) - 32 {IntDivResultM[31]}}, IntDivResultM[31:0]}),
					.s(W64M),
					.y(FIntDivResultM)
				);
			end
			else begin : genblk1
				assign FIntDivResultM = IntDivResultM[$signed(P[4216-:32]) - 1:0];
			end
		end
		else begin : genblk2
			assign FIntDivResultM = 1'sb0;
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module fdivsqrtpreproc (
	clk,
	IFDivStartE,
	Xm,
	Ym,
	Xe,
	Ye,
	FmtE,
	Bias,
	Nf,
	SqrtE,
	XZeroE,
	Funct3E,
	UeM,
	X,
	D,
	ForwardedSrcAE,
	ForwardedSrcBE,
	IntDivE,
	W64E,
	ISpecialCaseE,
	CyclesE,
	IntNormShiftM,
	ALTBM,
	W64M,
	AsM,
	BsM,
	BZeroM,
	AM
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire IFDivStartE;
	input wire [$signed(P[805-:32]):0] Xm;
	input wire [$signed(P[805-:32]):0] Ym;
	input wire [$signed(P[837-:32]) - 1:0] Xe;
	input wire [$signed(P[837-:32]) - 1:0] Ye;
	input wire [$signed(P[707-:32]) - 1:0] FmtE;
	input wire [$signed(P[837-:32]) - 2:0] Bias;
	input wire [$signed(P[869-:32]) - 1:0] Nf;
	input wire SqrtE;
	input wire XZeroE;
	input wire [2:0] Funct3E;
	output wire [$signed(P[837-:32]) + 1:0] UeM;
	output wire [$signed(P[95-:32]) + 3:0] X;
	output wire [$signed(P[95-:32]) + 3:0] D;
	input wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcAE;
	input wire [$signed(P[4216-:32]) - 1:0] ForwardedSrcBE;
	input wire IntDivE;
	input wire W64E;
	output wire ISpecialCaseE;
	output wire [$signed(P[127-:32]) - 1:0] CyclesE;
	output wire [$signed(P[63-:32]) - 1:0] IntNormShiftM;
	output wire ALTBM;
	output wire W64M;
	output wire AsM;
	output wire BsM;
	output wire BZeroM;
	output wire [$signed(P[4216-:32]) - 1:0] AM;
	wire [$signed(P[95-:32]):0] Xnorm;
	wire [$signed(P[95-:32]):0] Dnorm;
	wire [$signed(P[95-:32]) + 3:0] DivX;
	wire [$signed(P[95-:32]) + 3:0] DivXShifted;
	wire [$signed(P[95-:32]) + 3:0] SqrtX;
	wire [$signed(P[95-:32]) + 3:0] PreShiftX;
	wire [$signed(P[837-:32]) + 1:0] UeE;
	wire [$signed(P[95-:32]):0] IFX;
	wire [$signed(P[95-:32]):0] IFD;
	wire [$signed(P[63-:32]) - 1:0] mE;
	wire [$signed(P[63-:32]) - 1:0] ell;
	wire [$signed(P[63-:32]) - 1:0] IntResultBitsE;
	wire AZeroE;
	wire BZeroE;
	wire SignedDivE;
	wire AsE;
	wire BsE;
	wire [$signed(P[4216-:32]) - 1:0] AE;
	wire ALTBE;
	wire EvenExp;
	generate
		if (P[3729]) begin : intpreproc
			wire [$signed(P[4216-:32]) - 1:0] BE;
			wire [$signed(P[4216-:32]) - 1:0] PosA;
			wire [$signed(P[4216-:32]) - 1:0] PosB;
			assign SignedDivE = ~Funct3E[0];
			if ($signed(P[4216-:32]) == 64) begin : genblk1
				mux2 #(.WIDTH(64)) amux(
					.d0(ForwardedSrcAE),
					.d1({{32 {ForwardedSrcAE[31] & SignedDivE}}, ForwardedSrcAE[31:0]}),
					.s(W64E),
					.y(AE)
				);
				mux2 #(.WIDTH(64)) bmux(
					.d0(ForwardedSrcBE),
					.d1({{32 {ForwardedSrcBE[31] & SignedDivE}}, ForwardedSrcBE[31:0]}),
					.s(W64E),
					.y(BE)
				);
			end
			else begin : genblk1
				assign AE = ForwardedSrcAE;
				assign BE = ForwardedSrcBE;
			end
			assign AZeroE = ~(|AE);
			assign BZeroE = ~(|BE);
			assign AsE = AE[$signed(P[4216-:32]) - 1] & SignedDivE;
			assign BsE = BE[$signed(P[4216-:32]) - 1] & SignedDivE;
			mux2 #(.WIDTH($signed(P[4216-:32]))) posamux(
				.d0(AE),
				.d1(-AE),
				.s(AsE),
				.y(PosA)
			);
			mux2 #(.WIDTH($signed(P[4216-:32]))) posbmux(
				.d0(BE),
				.d1(-BE),
				.s(BsE),
				.y(PosB)
			);
			mux2 #(.WIDTH($signed(P[95-:32]) + 1)) ifxmux(
				.d0({Xm, {$signed(P[95-:32]) - $signed(P[805-:32]) {1'b0}}}),
				.d1({PosA, {($signed(P[95-:32]) - $signed(P[4216-:32])) + 1 {1'b0}}}),
				.s(IntDivE),
				.y(IFX)
			);
			mux2 #(.WIDTH($signed(P[95-:32]) + 1)) ifdmux(
				.d0({Ym, {$signed(P[95-:32]) - $signed(P[805-:32]) {1'b0}}}),
				.d1({PosB, {($signed(P[95-:32]) - $signed(P[4216-:32])) + 1 {1'b0}}}),
				.s(IntDivE),
				.y(IFD)
			);
		end
		else begin : genblk1
			assign IFX = {Xm, {$signed(P[95-:32]) - $signed(P[805-:32]) {1'b0}}};
			assign IFD = {Ym, {$signed(P[95-:32]) - $signed(P[805-:32]) {1'b0}}};
		end
	endgenerate
	lzc #(.WIDTH($signed(P[95-:32]) + 1)) lzcX(
		.num(IFX),
		.ZeroCnt(ell)
	);
	lzc #(.WIDTH($signed(P[95-:32]) + 1)) lzcY(
		.num(IFD),
		.ZeroCnt(mE)
	);
	assign Xnorm = IFX << ell;
	assign Dnorm = IFD << mE;
	generate
		if (P[3729]) begin : intrightshift
			wire [$signed(P[63-:32]) - 1:0] ZeroDiff;
			wire [$signed(P[63-:32]) - 1:0] p;
			assign ZeroDiff = mE - ell;
			assign ALTBE = ZeroDiff[$signed(P[63-:32]) - 1];
			localparam sv2v_uu_pmux_WIDTH = $signed(P[63-:32]);
			localparam [sv2v_uu_pmux_WIDTH - 1:0] sv2v_uu_pmux_ext_d1_0 = 1'sb0;
			mux2 #(.WIDTH($signed(P[63-:32]))) pmux(
				.d0(ZeroDiff),
				.d1(sv2v_uu_pmux_ext_d1_0),
				.s(ALTBE),
				.y(p)
			);
			assign IntResultBitsE = $signed(P[223-:32]) + p;
			assign ISpecialCaseE = BZeroE | ALTBE;
			if ($signed(P[191-:32]) > 1) begin : genblk1
				wire [$clog2($signed(P[191-:32])) - 1:0] RightShiftX;
				assign RightShiftX = ($signed(P[191-:32]) - 1) - ((IntResultBitsE - 1) % $signed(P[191-:32]));
				assign DivXShifted = DivX >> RightShiftX;
			end
			else begin : genblk1
				assign DivXShifted = DivX;
			end
		end
		else begin : genblk2
			assign {ISpecialCaseE, IntResultBitsE} = 1'sb0;
		end
	endgenerate
	assign DivX = {3'b000, Xnorm};
	assign EvenExp = Xe[0] ^ ell[0];
	mux2 #(.WIDTH($signed(P[95-:32]) + 4)) sqrtxmux(
		.d0({4'b0000, Xnorm[$signed(P[95-:32]):1]}),
		.d1({5'b00000, Xnorm[$signed(P[95-:32]):2]}),
		.s(EvenExp),
		.y(SqrtX)
	);
	mux2 #(.WIDTH($signed(P[95-:32]) + 4)) prexmux(
		.d0(DivX),
		.d1(SqrtX),
		.s(SqrtE),
		.y(PreShiftX)
	);
	generate
		if (P[3729]) begin : genblk3
			mux2 #(.WIDTH($signed(P[95-:32]) + 4)) xmux(
				.d0(PreShiftX),
				.d1(DivXShifted),
				.s(IntDivE),
				.y(X)
			);
		end
		else begin : genblk3
			assign X = PreShiftX;
		end
	endgenerate
	flopen #(.WIDTH($signed(P[95-:32]) + 4)) dreg(
		.clk(clk),
		.en(IFDivStartE),
		.d({3'b000, Dnorm}),
		.q(D)
	);
	fdivsqrtexpcalc #(.P(P)) expcalc(
		.Bias(Bias),
		.Xe(Xe),
		.Ye(Ye),
		.Sqrt(SqrtE),
		.ell(ell),
		.m(mE),
		.Ue(UeE)
	);
	flopen #(.WIDTH($signed(P[837-:32]) + 2)) expreg(
		.clk(clk),
		.en(IFDivStartE),
		.d(UeE),
		.q(UeM)
	);
	fdivsqrtcycles #(.P(P)) cyclecalc(
		.Nf(Nf),
		.IntDivE(IntDivE),
		.IntResultBitsE(IntResultBitsE),
		.CyclesE(CyclesE)
	);
	generate
		if (P[3729]) begin : intpipelineregs
			wire [$signed(P[63-:32]) - 1:0] IntDivNormShiftE;
			wire [$signed(P[63-:32]) - 1:0] IntRemNormShiftE;
			wire [$signed(P[63-:32]) - 1:0] IntNormShiftE;
			wire RemOpE;
			assign IntDivNormShiftE = $signed(P[31-:32]) - ((CyclesE * $signed(P[191-:32])) - $signed(P[223-:32]));
			assign IntRemNormShiftE = mE + ($signed(P[31-:32]) - ($signed(P[4216-:32]) - 1));
			assign RemOpE = Funct3E[1];
			mux2 #(.WIDTH($signed(P[63-:32]))) normshiftmux(
				.d0(IntDivNormShiftE),
				.d1(IntRemNormShiftE),
				.s(RemOpE),
				.y(IntNormShiftE)
			);
			flopen #(.WIDTH(1)) altbreg(
				.clk(clk),
				.en(IFDivStartE),
				.d(ALTBE),
				.q(ALTBM)
			);
			flopen #(.WIDTH(1)) bzeroreg(
				.clk(clk),
				.en(IFDivStartE),
				.d(BZeroE),
				.q(BZeroM)
			);
			flopen #(.WIDTH(1)) asignreg(
				.clk(clk),
				.en(IFDivStartE),
				.d(AsE),
				.q(AsM)
			);
			flopen #(.WIDTH(1)) bsignreg(
				.clk(clk),
				.en(IFDivStartE),
				.d(BsE),
				.q(BsM)
			);
			flopen #(.WIDTH($signed(P[63-:32]))) nsreg(
				.clk(clk),
				.en(IFDivStartE),
				.d(IntNormShiftE),
				.q(IntNormShiftM)
			);
			flopen #(.WIDTH($signed(P[4216-:32]))) srcareg(
				.clk(clk),
				.en(IFDivStartE),
				.d(AE),
				.q(AM)
			);
			if ($signed(P[4216-:32]) == 64) begin : genblk1
				flopen #(.WIDTH(1)) w64reg(
					.clk(clk),
					.en(IFDivStartE),
					.d(W64E),
					.q(W64M)
				);
			end
			else begin : genblk1
				assign W64M = 0;
			end
		end
		else begin : genblk4
			assign {ALTBM, W64M, AsM, BsM, BZeroM, AM, IntNormShiftM} = 1'sb0;
		end
	endgenerate
endmodule
module fdivsqrtstage2 (
	D,
	DBar,
	U,
	UM,
	WS,
	WC,
	C,
	SqrtE,
	un,
	CNext,
	UNext,
	UMNext,
	WSNext,
	WCNext
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[95-:32]) + 3:0] D;
	input wire [$signed(P[95-:32]) + 3:0] DBar;
	input wire [$signed(P[95-:32]):0] U;
	input wire [$signed(P[95-:32]):0] UM;
	input wire [$signed(P[95-:32]) + 3:0] WS;
	input wire [$signed(P[95-:32]) + 3:0] WC;
	input wire [$signed(P[95-:32]) + 1:0] C;
	input wire SqrtE;
	output wire un;
	output wire [$signed(P[95-:32]) + 1:0] CNext;
	output wire [$signed(P[95-:32]):0] UNext;
	output wire [$signed(P[95-:32]):0] UMNext;
	output wire [$signed(P[95-:32]) + 3:0] WSNext;
	output wire [$signed(P[95-:32]) + 3:0] WCNext;
	reg [$signed(P[95-:32]) + 3:0] Dsel;
	wire up;
	wire uz;
	wire [$signed(P[95-:32]) + 3:0] F;
	wire [$signed(P[95-:32]) + 3:0] AddIn;
	wire [$signed(P[95-:32]) + 3:0] WSA;
	wire [$signed(P[95-:32]) + 3:0] WCA;
	fdivsqrtuslc2 uslc2(
		.WS(WS[$signed(P[95-:32]) + 3:$signed(P[95-:32])]),
		.WC(WC[$signed(P[95-:32]) + 3:$signed(P[95-:32])]),
		.up(up),
		.uz(uz),
		.un(un)
	);
	fdivsqrtfgen2 #(.P(P)) fgen2(
		.up(up),
		.uz(uz),
		.C({2'b11, CNext}),
		.U({3'b000, U}),
		.UM({3'b000, UM}),
		.F(F)
	);
	always @(*) begin
		if (_sv2v_0)
			;
		if (up)
			Dsel = DBar;
		else if (uz)
			Dsel = 1'sb0;
		else
			Dsel = D;
	end
	mux2 #(.WIDTH($signed(P[95-:32]) + 4)) addinmux(
		.d0(Dsel),
		.d1(F),
		.s(SqrtE),
		.y(AddIn)
	);
	csa #(.N($signed(P[95-:32]) + 4)) csa(
		.x(WS),
		.y(WC),
		.z(AddIn),
		.cin(up & ~SqrtE),
		.s(WSA),
		.c(WCA)
	);
	assign WSNext = WSA << 1;
	assign WCNext = WCA << 1;
	assign CNext = {1'b1, C[$signed(P[95-:32]) + 1:1]};
	fdivsqrtuotfc2 #(.P(P)) uotfc2(
		.up(up),
		.un(un),
		.C(CNext),
		.U(U),
		.UM(UM),
		.UNext(UNext),
		.UMNext(UMNext)
	);
	initial _sv2v_0 = 0;
endmodule
module fdivsqrtstage4 (
	D,
	DBar,
	D2,
	DBar2,
	U,
	UM,
	WS,
	WC,
	C,
	SqrtE,
	CNext,
	un,
	UNext,
	UMNext,
	WSNext,
	WCNext
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[95-:32]) + 3:0] D;
	input wire [$signed(P[95-:32]) + 3:0] DBar;
	input wire [$signed(P[95-:32]) + 3:0] D2;
	input wire [$signed(P[95-:32]) + 3:0] DBar2;
	input wire [$signed(P[95-:32]):0] U;
	input wire [$signed(P[95-:32]):0] UM;
	input wire [$signed(P[95-:32]) + 3:0] WS;
	input wire [$signed(P[95-:32]) + 3:0] WC;
	input wire [$signed(P[95-:32]) + 1:0] C;
	input wire SqrtE;
	output wire [$signed(P[95-:32]) + 1:0] CNext;
	output wire un;
	output wire [$signed(P[95-:32]):0] UNext;
	output wire [$signed(P[95-:32]):0] UMNext;
	output wire [$signed(P[95-:32]) + 3:0] WSNext;
	output wire [$signed(P[95-:32]) + 3:0] WCNext;
	reg [$signed(P[95-:32]) + 3:0] Dsel;
	wire [3:0] udigit;
	wire [$signed(P[95-:32]) + 3:0] F;
	wire [$signed(P[95-:32]) + 3:0] AddIn;
	wire [4:0] Smsbs;
	wire [2:0] Dmsbs;
	wire [7:0] WCmsbs;
	wire [7:0] WSmsbs;
	wire CarryIn;
	wire [$signed(P[95-:32]) + 3:0] WSA;
	wire [$signed(P[95-:32]) + 3:0] WCA;
	wire j0;
	wire j1;
	assign j0 = ~C[$signed(P[95-:32]) + 1];
	assign j1 = ~C[$signed(P[95-:32]) - 1];
	assign Smsbs = U[$signed(P[95-:32]):$signed(P[95-:32]) - 4];
	assign Dmsbs = D[$signed(P[95-:32]) - 1:$signed(P[95-:32]) - 3];
	assign WCmsbs = WC[$signed(P[95-:32]) + 3:$signed(P[95-:32]) - 4];
	assign WSmsbs = WS[$signed(P[95-:32]) + 3:$signed(P[95-:32]) - 4];
	fdivsqrtuslc4cmp uslc4(
		.Dmsbs(Dmsbs),
		.Smsbs(Smsbs),
		.WSmsbs(WSmsbs),
		.WCmsbs(WCmsbs),
		.SqrtE(SqrtE),
		.j0(j0),
		.j1(j1),
		.udigit(udigit)
	);
	assign un = 1'b0;
	fdivsqrtfgen4 #(.P(P)) fgen4(
		.udigit(udigit),
		.C({2'b11, CNext}),
		.U({3'b000, U}),
		.UM({3'b000, UM}),
		.F(F)
	);
	always @(*) begin
		if (_sv2v_0)
			;
		case (udigit)
			4'b1000: Dsel = DBar2;
			4'b0100: Dsel = DBar;
			4'b0000: Dsel = 1'sb0;
			4'b0010: Dsel = D;
			4'b0001: Dsel = D2;
			default: Dsel = 1'sbx;
		endcase
	end
	assign AddIn = (SqrtE ? F : Dsel);
	assign CarryIn = ~SqrtE & (udigit[3] | udigit[2]);
	csa #(.N($signed(P[95-:32]) + 4)) csa(
		.x(WS),
		.y(WC),
		.z(AddIn),
		.cin(CarryIn),
		.s(WSA),
		.c(WCA)
	);
	assign WSNext = WSA << 2;
	assign WCNext = WCA << 2;
	assign CNext = {2'b11, C[$signed(P[95-:32]) + 1:2]};
	fdivsqrtuotfc4 #(.P(P)) fdivsqrtuotfc4(
		.udigit(udigit),
		.C(CNext[$signed(P[95-:32]):0]),
		.U(U),
		.UM(UM),
		.UNext(UNext),
		.UMNext(UMNext)
	);
	initial _sv2v_0 = 0;
endmodule
module fdivsqrtuotfc2 (
	up,
	un,
	C,
	U,
	UM,
	UNext,
	UMNext
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire up;
	input wire un;
	input wire [$signed(P[95-:32]) + 1:0] C;
	input wire [$signed(P[95-:32]):0] U;
	input wire [$signed(P[95-:32]):0] UM;
	output reg [$signed(P[95-:32]):0] UNext;
	output reg [$signed(P[95-:32]):0] UMNext;
	wire [$signed(P[95-:32]):0] K;
	assign K = C[$signed(P[95-:32]):0] & ~(C[$signed(P[95-:32]):0] << 1);
	always @(*) begin
		if (_sv2v_0)
			;
		if (up) begin
			UNext = U | K;
			UMNext = U;
		end
		else if (un) begin
			UNext = UM | K;
			UMNext = UM;
		end
		else begin
			UNext = U;
			UMNext = UM | K;
		end
	end
	initial _sv2v_0 = 0;
endmodule
module fdivsqrtuotfc4 (
	udigit,
	U,
	UM,
	C,
	UNext,
	UMNext
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [3:0] udigit;
	input wire [$signed(P[95-:32]):0] U;
	input wire [$signed(P[95-:32]):0] UM;
	input wire [$signed(P[95-:32]):0] C;
	output reg [$signed(P[95-:32]):0] UNext;
	output reg [$signed(P[95-:32]):0] UMNext;
	wire [$signed(P[95-:32]):0] K1;
	wire [$signed(P[95-:32]):0] K2;
	wire [$signed(P[95-:32]):0] K3;
	assign K1 = C & ~(C << 1);
	assign K2 = (C << 1) & ~(C << 2);
	assign K3 = C & ~(C << 2);
	always @(*) begin
		if (_sv2v_0)
			;
		if (udigit[3]) begin
			UNext = U | K2;
			UMNext = U | K1;
		end
		else if (udigit[2]) begin
			UNext = U | K1;
			UMNext = U;
		end
		else if (udigit[1]) begin
			UNext = UM | K3;
			UMNext = UM | K2;
		end
		else if (udigit[0]) begin
			UNext = UM | K2;
			UMNext = UM | K1;
		end
		else begin
			UNext = U;
			UMNext = UM | K3;
		end
	end
	initial _sv2v_0 = 0;
endmodule
module fdivsqrtuslc2 (
	WS,
	WC,
	up,
	uz,
	un
);
	input wire [3:0] WS;
	input wire [3:0] WC;
	output wire up;
	output wire uz;
	output wire un;
	wire sign;
	assign uz = ((WS[2] ^ WC[2]) & (WS[1] ^ WC[1])) & (WS[0] ^ WC[0]);
	assign sign = (WS[3] ^ WC[3]) ^ ((WS[2] & WC[2]) | ((WS[2] ^ WC[2]) & ((WS[1] & WC[1]) | ((WS[1] ^ WC[1]) & (WS[0] & WC[0])))));
	assign up = ~uz & ~sign;
	assign un = ~uz & sign;
endmodule
module fdivsqrtuslc4cmp (
	Dmsbs,
	Smsbs,
	WSmsbs,
	WCmsbs,
	SqrtE,
	j0,
	j1,
	udigit
);
	reg _sv2v_0;
	input wire [2:0] Dmsbs;
	input wire [4:0] Smsbs;
	input wire [7:0] WSmsbs;
	input wire [7:0] WCmsbs;
	input wire SqrtE;
	input wire j0;
	input wire j1;
	output reg [3:0] udigit;
	wire [6:0] Wmsbs;
	wire [7:0] PreWmsbs;
	reg [2:0] A;
	assign PreWmsbs = WCmsbs + WSmsbs;
	assign Wmsbs = PreWmsbs[7:1];
	wire [6:0] mk2;
	wire [6:0] mk1;
	wire [6:0] mk0;
	wire [6:0] mkm1;
	wire [6:0] mkj2;
	wire [6:0] mkj1;
	wire [6:0] mks2 [7:0];
	wire [6:0] mks1 [7:0];
	wire [6:0] mks0 [7:0];
	wire [6:0] mksm1 [7:0];
	wire sqrtspecial;
	assign mks2[0] = 12;
	assign mks2[1] = 14;
	assign mks2[2] = 16;
	assign mks2[3] = 17;
	assign mks2[4] = 18;
	assign mks2[5] = 20;
	assign mks2[6] = 22;
	assign mks2[7] = 23;
	assign mks1[0] = 4;
	assign mks1[1] = 4;
	assign mks1[2] = 6;
	assign mks1[3] = 6;
	assign mks1[4] = 6;
	assign mks1[5] = 8;
	assign mks1[6] = 8;
	assign mks1[7] = 8;
	assign mks0[0] = -4;
	assign mks0[1] = -4;
	assign mks0[2] = -6;
	assign mks0[3] = -6;
	assign mks0[4] = -6;
	assign mks0[5] = -8;
	assign mks0[6] = -8;
	assign mks0[7] = -8;
	assign mksm1[0] = -13;
	assign mksm1[1] = -14;
	assign mksm1[2] = -16;
	assign mksm1[3] = -17;
	assign mksm1[4] = -18;
	assign mksm1[5] = -20;
	assign mksm1[6] = -22;
	assign mksm1[7] = -23;
	assign mkj2 = 20;
	assign mkj1 = (j0 ? 0 : 8);
	assign sqrtspecial = SqrtE & (j1 | j0);
	always @(*) begin
		if (_sv2v_0)
			;
		if (SqrtE) begin
			if (Smsbs[4])
				A = 3'b111;
			else
				A = Smsbs[2:0];
		end
		else
			A = Dmsbs;
	end
	assign mk2 = (sqrtspecial ? mkj2 : mks2[A]);
	assign mk1 = (sqrtspecial ? mkj1 : mks1[A]);
	assign mk0 = (sqrtspecial ? -mkj1 : mks0[A]);
	assign mkm1 = (sqrtspecial ? -mkj2 : mksm1[A]);
	always @(*) begin
		if (_sv2v_0)
			;
		if ($signed(Wmsbs) >= $signed(mk2))
			udigit = 4'b1000;
		else if ($signed(Wmsbs) >= $signed(mk1))
			udigit = 4'b0100;
		else if ($signed(Wmsbs) >= $signed(mk0))
			udigit = 4'b0000;
		else if ($signed(Wmsbs) >= $signed(mkm1))
			udigit = 4'b0010;
		else
			udigit = 4'b0001;
	end
	initial _sv2v_0 = 0;
endmodule
module fdivsqrtuslc4 (
	Dmsbs,
	Smsbs,
	WSmsbs,
	WCmsbs,
	Sqrt,
	j0,
	j1,
	udigit
);
	reg _sv2v_0;
	input wire [2:0] Dmsbs;
	input wire [4:0] Smsbs;
	input wire [7:0] WSmsbs;
	input wire [7:0] WCmsbs;
	input wire Sqrt;
	input wire j0;
	input wire j1;
	output wire [3:0] udigit;
	wire [7:0] PreWmsbs;
	wire [6:0] Wmsbs;
	reg [2:0] A;
	assign PreWmsbs = WCmsbs + WSmsbs;
	assign Wmsbs = PreWmsbs[7:1];
	reg [3:0] USel4;
	always @(*) begin : sv2v_autoblock_1
		case ({A, Wmsbs})
			10'd0: USel4 = 4'b0000;
			10'd1: USel4 = 4'b0000;
			10'd2: USel4 = 4'b0000;
			10'd3: USel4 = 4'b0000;
			10'd4: USel4 = 4'b0100;
			10'd5: USel4 = 4'b0100;
			10'd6: USel4 = 4'b0100;
			10'd7: USel4 = 4'b0100;
			10'd8: USel4 = 4'b0100;
			10'd9: USel4 = 4'b0100;
			10'd10: USel4 = 4'b0100;
			10'd11: USel4 = 4'b0100;
			10'd12: USel4 = 4'b1000;
			10'd13: USel4 = 4'b1000;
			10'd14: USel4 = 4'b1000;
			10'd15: USel4 = 4'b1000;
			10'd16: USel4 = 4'b1000;
			10'd17: USel4 = 4'b1000;
			10'd18: USel4 = 4'b1000;
			10'd19: USel4 = 4'b1000;
			10'd20: USel4 = 4'b1000;
			10'd21: USel4 = 4'b1000;
			10'd22: USel4 = 4'b1000;
			10'd23: USel4 = 4'b1000;
			10'd24: USel4 = 4'b1000;
			10'd25: USel4 = 4'b1000;
			10'd26: USel4 = 4'b1000;
			10'd27: USel4 = 4'b1000;
			10'd28: USel4 = 4'b1000;
			10'd29: USel4 = 4'b1000;
			10'd30: USel4 = 4'b1000;
			10'd31: USel4 = 4'b1000;
			10'd32: USel4 = 4'b1000;
			10'd33: USel4 = 4'b1000;
			10'd34: USel4 = 4'b1000;
			10'd35: USel4 = 4'b1000;
			10'd36: USel4 = 4'b1000;
			10'd37: USel4 = 4'b1000;
			10'd38: USel4 = 4'b1000;
			10'd39: USel4 = 4'b1000;
			10'd40: USel4 = 4'b1000;
			10'd41: USel4 = 4'b1000;
			10'd42: USel4 = 4'b1000;
			10'd43: USel4 = 4'b1000;
			10'd44: USel4 = 4'b1000;
			10'd45: USel4 = 4'b1000;
			10'd46: USel4 = 4'b1000;
			10'd47: USel4 = 4'b1000;
			10'd48: USel4 = 4'b1000;
			10'd49: USel4 = 4'b1000;
			10'd50: USel4 = 4'b1000;
			10'd51: USel4 = 4'b1000;
			10'd52: USel4 = 4'b1000;
			10'd53: USel4 = 4'b1000;
			10'd54: USel4 = 4'b1000;
			10'd55: USel4 = 4'b1000;
			10'd56: USel4 = 4'b1000;
			10'd57: USel4 = 4'b1000;
			10'd58: USel4 = 4'b1000;
			10'd59: USel4 = 4'b1000;
			10'd60: USel4 = 4'b1000;
			10'd61: USel4 = 4'b1000;
			10'd62: USel4 = 4'b1000;
			10'd63: USel4 = 4'b1000;
			10'd64: USel4 = 4'b0001;
			10'd65: USel4 = 4'b0001;
			10'd66: USel4 = 4'b0001;
			10'd67: USel4 = 4'b0001;
			10'd68: USel4 = 4'b0001;
			10'd69: USel4 = 4'b0001;
			10'd70: USel4 = 4'b0001;
			10'd71: USel4 = 4'b0001;
			10'd72: USel4 = 4'b0001;
			10'd73: USel4 = 4'b0001;
			10'd74: USel4 = 4'b0001;
			10'd75: USel4 = 4'b0001;
			10'd76: USel4 = 4'b0001;
			10'd77: USel4 = 4'b0001;
			10'd78: USel4 = 4'b0001;
			10'd79: USel4 = 4'b0001;
			10'd80: USel4 = 4'b0001;
			10'd81: USel4 = 4'b0001;
			10'd82: USel4 = 4'b0001;
			10'd83: USel4 = 4'b0001;
			10'd84: USel4 = 4'b0001;
			10'd85: USel4 = 4'b0001;
			10'd86: USel4 = 4'b0001;
			10'd87: USel4 = 4'b0001;
			10'd88: USel4 = 4'b0001;
			10'd89: USel4 = 4'b0001;
			10'd90: USel4 = 4'b0001;
			10'd91: USel4 = 4'b0001;
			10'd92: USel4 = 4'b0001;
			10'd93: USel4 = 4'b0001;
			10'd94: USel4 = 4'b0001;
			10'd95: USel4 = 4'b0001;
			10'd96: USel4 = 4'b0001;
			10'd97: USel4 = 4'b0001;
			10'd98: USel4 = 4'b0001;
			10'd99: USel4 = 4'b0001;
			10'd100: USel4 = 4'b0001;
			10'd101: USel4 = 4'b0001;
			10'd102: USel4 = 4'b0001;
			10'd103: USel4 = 4'b0001;
			10'd104: USel4 = 4'b0001;
			10'd105: USel4 = 4'b0001;
			10'd106: USel4 = 4'b0001;
			10'd107: USel4 = 4'b0001;
			10'd108: USel4 = 4'b0001;
			10'd109: USel4 = 4'b0001;
			10'd110: USel4 = 4'b0001;
			10'd111: USel4 = 4'b0001;
			10'd112: USel4 = 4'b0001;
			10'd113: USel4 = 4'b0001;
			10'd114: USel4 = 4'b0001;
			10'd115: USel4 = 4'b0010;
			10'd116: USel4 = 4'b0010;
			10'd117: USel4 = 4'b0010;
			10'd118: USel4 = 4'b0010;
			10'd119: USel4 = 4'b0010;
			10'd120: USel4 = 4'b0010;
			10'd121: USel4 = 4'b0010;
			10'd122: USel4 = 4'b0010;
			10'd123: USel4 = 4'b0010;
			10'd124: USel4 = 4'b0000;
			10'd125: USel4 = 4'b0000;
			10'd126: USel4 = 4'b0000;
			10'd127: USel4 = 4'b0000;
			10'd128: USel4 = 4'b0000;
			10'd129: USel4 = 4'b0000;
			10'd130: USel4 = 4'b0000;
			10'd131: USel4 = 4'b0000;
			10'd132: USel4 = 4'b0100;
			10'd133: USel4 = 4'b0100;
			10'd134: USel4 = 4'b0100;
			10'd135: USel4 = 4'b0100;
			10'd136: USel4 = 4'b0100;
			10'd137: USel4 = 4'b0100;
			10'd138: USel4 = 4'b0100;
			10'd139: USel4 = 4'b0100;
			10'd140: USel4 = 4'b0100;
			10'd141: USel4 = 4'b0100;
			10'd142: USel4 = 4'b1000;
			10'd143: USel4 = 4'b1000;
			10'd144: USel4 = 4'b1000;
			10'd145: USel4 = 4'b1000;
			10'd146: USel4 = 4'b1000;
			10'd147: USel4 = 4'b1000;
			10'd148: USel4 = 4'b1000;
			10'd149: USel4 = 4'b1000;
			10'd150: USel4 = 4'b1000;
			10'd151: USel4 = 4'b1000;
			10'd152: USel4 = 4'b1000;
			10'd153: USel4 = 4'b1000;
			10'd154: USel4 = 4'b1000;
			10'd155: USel4 = 4'b1000;
			10'd156: USel4 = 4'b1000;
			10'd157: USel4 = 4'b1000;
			10'd158: USel4 = 4'b1000;
			10'd159: USel4 = 4'b1000;
			10'd160: USel4 = 4'b1000;
			10'd161: USel4 = 4'b1000;
			10'd162: USel4 = 4'b1000;
			10'd163: USel4 = 4'b1000;
			10'd164: USel4 = 4'b1000;
			10'd165: USel4 = 4'b1000;
			10'd166: USel4 = 4'b1000;
			10'd167: USel4 = 4'b1000;
			10'd168: USel4 = 4'b1000;
			10'd169: USel4 = 4'b1000;
			10'd170: USel4 = 4'b1000;
			10'd171: USel4 = 4'b1000;
			10'd172: USel4 = 4'b1000;
			10'd173: USel4 = 4'b1000;
			10'd174: USel4 = 4'b1000;
			10'd175: USel4 = 4'b1000;
			10'd176: USel4 = 4'b1000;
			10'd177: USel4 = 4'b1000;
			10'd178: USel4 = 4'b1000;
			10'd179: USel4 = 4'b1000;
			10'd180: USel4 = 4'b1000;
			10'd181: USel4 = 4'b1000;
			10'd182: USel4 = 4'b1000;
			10'd183: USel4 = 4'b1000;
			10'd184: USel4 = 4'b1000;
			10'd185: USel4 = 4'b1000;
			10'd186: USel4 = 4'b1000;
			10'd187: USel4 = 4'b1000;
			10'd188: USel4 = 4'b1000;
			10'd189: USel4 = 4'b1000;
			10'd190: USel4 = 4'b1000;
			10'd191: USel4 = 4'b1000;
			10'd192: USel4 = 4'b0001;
			10'd193: USel4 = 4'b0001;
			10'd194: USel4 = 4'b0001;
			10'd195: USel4 = 4'b0001;
			10'd196: USel4 = 4'b0001;
			10'd197: USel4 = 4'b0001;
			10'd198: USel4 = 4'b0001;
			10'd199: USel4 = 4'b0001;
			10'd200: USel4 = 4'b0001;
			10'd201: USel4 = 4'b0001;
			10'd202: USel4 = 4'b0001;
			10'd203: USel4 = 4'b0001;
			10'd204: USel4 = 4'b0001;
			10'd205: USel4 = 4'b0001;
			10'd206: USel4 = 4'b0001;
			10'd207: USel4 = 4'b0001;
			10'd208: USel4 = 4'b0001;
			10'd209: USel4 = 4'b0001;
			10'd210: USel4 = 4'b0001;
			10'd211: USel4 = 4'b0001;
			10'd212: USel4 = 4'b0001;
			10'd213: USel4 = 4'b0001;
			10'd214: USel4 = 4'b0001;
			10'd215: USel4 = 4'b0001;
			10'd216: USel4 = 4'b0001;
			10'd217: USel4 = 4'b0001;
			10'd218: USel4 = 4'b0001;
			10'd219: USel4 = 4'b0001;
			10'd220: USel4 = 4'b0001;
			10'd221: USel4 = 4'b0001;
			10'd222: USel4 = 4'b0001;
			10'd223: USel4 = 4'b0001;
			10'd224: USel4 = 4'b0001;
			10'd225: USel4 = 4'b0001;
			10'd226: USel4 = 4'b0001;
			10'd227: USel4 = 4'b0001;
			10'd228: USel4 = 4'b0001;
			10'd229: USel4 = 4'b0001;
			10'd230: USel4 = 4'b0001;
			10'd231: USel4 = 4'b0001;
			10'd232: USel4 = 4'b0001;
			10'd233: USel4 = 4'b0001;
			10'd234: USel4 = 4'b0001;
			10'd235: USel4 = 4'b0001;
			10'd236: USel4 = 4'b0001;
			10'd237: USel4 = 4'b0001;
			10'd238: USel4 = 4'b0001;
			10'd239: USel4 = 4'b0001;
			10'd240: USel4 = 4'b0001;
			10'd241: USel4 = 4'b0001;
			10'd242: USel4 = 4'b0010;
			10'd243: USel4 = 4'b0010;
			10'd244: USel4 = 4'b0010;
			10'd245: USel4 = 4'b0010;
			10'd246: USel4 = 4'b0010;
			10'd247: USel4 = 4'b0010;
			10'd248: USel4 = 4'b0010;
			10'd249: USel4 = 4'b0010;
			10'd250: USel4 = 4'b0010;
			10'd251: USel4 = 4'b0010;
			10'd252: USel4 = 4'b0000;
			10'd253: USel4 = 4'b0000;
			10'd254: USel4 = 4'b0000;
			10'd255: USel4 = 4'b0000;
			10'd256: USel4 = 4'b0000;
			10'd257: USel4 = 4'b0000;
			10'd258: USel4 = 4'b0000;
			10'd259: USel4 = 4'b0000;
			10'd260: USel4 = 4'b0100;
			10'd261: USel4 = 4'b0100;
			10'd262: USel4 = 4'b0100;
			10'd263: USel4 = 4'b0100;
			10'd264: USel4 = 4'b0100;
			10'd265: USel4 = 4'b0100;
			10'd266: USel4 = 4'b0100;
			10'd267: USel4 = 4'b0100;
			10'd268: USel4 = 4'b0100;
			10'd269: USel4 = 4'b0100;
			10'd270: USel4 = 4'b0100;
			10'd271: USel4 = 4'b0100;
			10'd272: USel4 = 4'b1000;
			10'd273: USel4 = 4'b1000;
			10'd274: USel4 = 4'b1000;
			10'd275: USel4 = 4'b1000;
			10'd276: USel4 = 4'b1000;
			10'd277: USel4 = 4'b1000;
			10'd278: USel4 = 4'b1000;
			10'd279: USel4 = 4'b1000;
			10'd280: USel4 = 4'b1000;
			10'd281: USel4 = 4'b1000;
			10'd282: USel4 = 4'b1000;
			10'd283: USel4 = 4'b1000;
			10'd284: USel4 = 4'b1000;
			10'd285: USel4 = 4'b1000;
			10'd286: USel4 = 4'b1000;
			10'd287: USel4 = 4'b1000;
			10'd288: USel4 = 4'b1000;
			10'd289: USel4 = 4'b1000;
			10'd290: USel4 = 4'b1000;
			10'd291: USel4 = 4'b1000;
			10'd292: USel4 = 4'b1000;
			10'd293: USel4 = 4'b1000;
			10'd294: USel4 = 4'b1000;
			10'd295: USel4 = 4'b1000;
			10'd296: USel4 = 4'b1000;
			10'd297: USel4 = 4'b1000;
			10'd298: USel4 = 4'b1000;
			10'd299: USel4 = 4'b1000;
			10'd300: USel4 = 4'b1000;
			10'd301: USel4 = 4'b1000;
			10'd302: USel4 = 4'b1000;
			10'd303: USel4 = 4'b1000;
			10'd304: USel4 = 4'b1000;
			10'd305: USel4 = 4'b1000;
			10'd306: USel4 = 4'b1000;
			10'd307: USel4 = 4'b1000;
			10'd308: USel4 = 4'b1000;
			10'd309: USel4 = 4'b1000;
			10'd310: USel4 = 4'b1000;
			10'd311: USel4 = 4'b1000;
			10'd312: USel4 = 4'b1000;
			10'd313: USel4 = 4'b1000;
			10'd314: USel4 = 4'b1000;
			10'd315: USel4 = 4'b1000;
			10'd316: USel4 = 4'b1000;
			10'd317: USel4 = 4'b1000;
			10'd318: USel4 = 4'b1000;
			10'd319: USel4 = 4'b1000;
			10'd320: USel4 = 4'b0001;
			10'd321: USel4 = 4'b0001;
			10'd322: USel4 = 4'b0001;
			10'd323: USel4 = 4'b0001;
			10'd324: USel4 = 4'b0001;
			10'd325: USel4 = 4'b0001;
			10'd326: USel4 = 4'b0001;
			10'd327: USel4 = 4'b0001;
			10'd328: USel4 = 4'b0001;
			10'd329: USel4 = 4'b0001;
			10'd330: USel4 = 4'b0001;
			10'd331: USel4 = 4'b0001;
			10'd332: USel4 = 4'b0001;
			10'd333: USel4 = 4'b0001;
			10'd334: USel4 = 4'b0001;
			10'd335: USel4 = 4'b0001;
			10'd336: USel4 = 4'b0001;
			10'd337: USel4 = 4'b0001;
			10'd338: USel4 = 4'b0001;
			10'd339: USel4 = 4'b0001;
			10'd340: USel4 = 4'b0001;
			10'd341: USel4 = 4'b0001;
			10'd342: USel4 = 4'b0001;
			10'd343: USel4 = 4'b0001;
			10'd344: USel4 = 4'b0001;
			10'd345: USel4 = 4'b0001;
			10'd346: USel4 = 4'b0001;
			10'd347: USel4 = 4'b0001;
			10'd348: USel4 = 4'b0001;
			10'd349: USel4 = 4'b0001;
			10'd350: USel4 = 4'b0001;
			10'd351: USel4 = 4'b0001;
			10'd352: USel4 = 4'b0001;
			10'd353: USel4 = 4'b0001;
			10'd354: USel4 = 4'b0001;
			10'd355: USel4 = 4'b0001;
			10'd356: USel4 = 4'b0001;
			10'd357: USel4 = 4'b0001;
			10'd358: USel4 = 4'b0001;
			10'd359: USel4 = 4'b0001;
			10'd360: USel4 = 4'b0001;
			10'd361: USel4 = 4'b0001;
			10'd362: USel4 = 4'b0001;
			10'd363: USel4 = 4'b0001;
			10'd364: USel4 = 4'b0001;
			10'd365: USel4 = 4'b0001;
			10'd366: USel4 = 4'b0001;
			10'd367: USel4 = 4'b0001;
			10'd368: USel4 = 4'b0010;
			10'd369: USel4 = 4'b0010;
			10'd370: USel4 = 4'b0010;
			10'd371: USel4 = 4'b0010;
			10'd372: USel4 = 4'b0010;
			10'd373: USel4 = 4'b0010;
			10'd374: USel4 = 4'b0010;
			10'd375: USel4 = 4'b0010;
			10'd376: USel4 = 4'b0010;
			10'd377: USel4 = 4'b0010;
			10'd378: USel4 = 4'b0000;
			10'd379: USel4 = 4'b0000;
			10'd380: USel4 = 4'b0000;
			10'd381: USel4 = 4'b0000;
			10'd382: USel4 = 4'b0000;
			10'd383: USel4 = 4'b0000;
			10'd384: USel4 = 4'b0000;
			10'd385: USel4 = 4'b0000;
			10'd386: USel4 = 4'b0000;
			10'd387: USel4 = 4'b0000;
			10'd388: USel4 = 4'b0100;
			10'd389: USel4 = 4'b0100;
			10'd390: USel4 = 4'b0100;
			10'd391: USel4 = 4'b0100;
			10'd392: USel4 = 4'b0100;
			10'd393: USel4 = 4'b0100;
			10'd394: USel4 = 4'b0100;
			10'd395: USel4 = 4'b0100;
			10'd396: USel4 = 4'b0100;
			10'd397: USel4 = 4'b0100;
			10'd398: USel4 = 4'b0100;
			10'd399: USel4 = 4'b0100;
			10'd400: USel4 = 4'b1000;
			10'd401: USel4 = 4'b1000;
			10'd402: USel4 = 4'b1000;
			10'd403: USel4 = 4'b1000;
			10'd404: USel4 = 4'b1000;
			10'd405: USel4 = 4'b1000;
			10'd406: USel4 = 4'b1000;
			10'd407: USel4 = 4'b1000;
			10'd408: USel4 = 4'b1000;
			10'd409: USel4 = 4'b1000;
			10'd410: USel4 = 4'b1000;
			10'd411: USel4 = 4'b1000;
			10'd412: USel4 = 4'b1000;
			10'd413: USel4 = 4'b1000;
			10'd414: USel4 = 4'b1000;
			10'd415: USel4 = 4'b1000;
			10'd416: USel4 = 4'b1000;
			10'd417: USel4 = 4'b1000;
			10'd418: USel4 = 4'b1000;
			10'd419: USel4 = 4'b1000;
			10'd420: USel4 = 4'b1000;
			10'd421: USel4 = 4'b1000;
			10'd422: USel4 = 4'b1000;
			10'd423: USel4 = 4'b1000;
			10'd424: USel4 = 4'b1000;
			10'd425: USel4 = 4'b1000;
			10'd426: USel4 = 4'b1000;
			10'd427: USel4 = 4'b1000;
			10'd428: USel4 = 4'b1000;
			10'd429: USel4 = 4'b1000;
			10'd430: USel4 = 4'b1000;
			10'd431: USel4 = 4'b1000;
			10'd432: USel4 = 4'b1000;
			10'd433: USel4 = 4'b1000;
			10'd434: USel4 = 4'b1000;
			10'd435: USel4 = 4'b1000;
			10'd436: USel4 = 4'b1000;
			10'd437: USel4 = 4'b1000;
			10'd438: USel4 = 4'b1000;
			10'd439: USel4 = 4'b1000;
			10'd440: USel4 = 4'b1000;
			10'd441: USel4 = 4'b1000;
			10'd442: USel4 = 4'b1000;
			10'd443: USel4 = 4'b1000;
			10'd444: USel4 = 4'b1000;
			10'd445: USel4 = 4'b1000;
			10'd446: USel4 = 4'b1000;
			10'd447: USel4 = 4'b1000;
			10'd448: USel4 = 4'b0001;
			10'd449: USel4 = 4'b0001;
			10'd450: USel4 = 4'b0001;
			10'd451: USel4 = 4'b0001;
			10'd452: USel4 = 4'b0001;
			10'd453: USel4 = 4'b0001;
			10'd454: USel4 = 4'b0001;
			10'd455: USel4 = 4'b0001;
			10'd456: USel4 = 4'b0001;
			10'd457: USel4 = 4'b0001;
			10'd458: USel4 = 4'b0001;
			10'd459: USel4 = 4'b0001;
			10'd460: USel4 = 4'b0001;
			10'd461: USel4 = 4'b0001;
			10'd462: USel4 = 4'b0001;
			10'd463: USel4 = 4'b0001;
			10'd464: USel4 = 4'b0001;
			10'd465: USel4 = 4'b0001;
			10'd466: USel4 = 4'b0001;
			10'd467: USel4 = 4'b0001;
			10'd468: USel4 = 4'b0001;
			10'd469: USel4 = 4'b0001;
			10'd470: USel4 = 4'b0001;
			10'd471: USel4 = 4'b0001;
			10'd472: USel4 = 4'b0001;
			10'd473: USel4 = 4'b0001;
			10'd474: USel4 = 4'b0001;
			10'd475: USel4 = 4'b0001;
			10'd476: USel4 = 4'b0001;
			10'd477: USel4 = 4'b0001;
			10'd478: USel4 = 4'b0001;
			10'd479: USel4 = 4'b0001;
			10'd480: USel4 = 4'b0001;
			10'd481: USel4 = 4'b0001;
			10'd482: USel4 = 4'b0001;
			10'd483: USel4 = 4'b0001;
			10'd484: USel4 = 4'b0001;
			10'd485: USel4 = 4'b0001;
			10'd486: USel4 = 4'b0001;
			10'd487: USel4 = 4'b0001;
			10'd488: USel4 = 4'b0001;
			10'd489: USel4 = 4'b0001;
			10'd490: USel4 = 4'b0001;
			10'd491: USel4 = 4'b0001;
			10'd492: USel4 = 4'b0001;
			10'd493: USel4 = 4'b0001;
			10'd494: USel4 = 4'b0001;
			10'd495: USel4 = 4'b0010;
			10'd496: USel4 = 4'b0010;
			10'd497: USel4 = 4'b0010;
			10'd498: USel4 = 4'b0010;
			10'd499: USel4 = 4'b0010;
			10'd500: USel4 = 4'b0010;
			10'd501: USel4 = 4'b0010;
			10'd502: USel4 = 4'b0010;
			10'd503: USel4 = 4'b0010;
			10'd504: USel4 = 4'b0010;
			10'd505: USel4 = 4'b0010;
			10'd506: USel4 = 4'b0000;
			10'd507: USel4 = 4'b0000;
			10'd508: USel4 = 4'b0000;
			10'd509: USel4 = 4'b0000;
			10'd510: USel4 = 4'b0000;
			10'd511: USel4 = 4'b0000;
			10'd512: USel4 = 4'b0000;
			10'd513: USel4 = 4'b0000;
			10'd514: USel4 = 4'b0000;
			10'd515: USel4 = 4'b0000;
			10'd516: USel4 = 4'b0000;
			10'd517: USel4 = 4'b0000;
			10'd518: USel4 = 4'b0100;
			10'd519: USel4 = 4'b0100;
			10'd520: USel4 = 4'b0100;
			10'd521: USel4 = 4'b0100;
			10'd522: USel4 = 4'b0100;
			10'd523: USel4 = 4'b0100;
			10'd524: USel4 = 4'b0100;
			10'd525: USel4 = 4'b0100;
			10'd526: USel4 = 4'b0100;
			10'd527: USel4 = 4'b0100;
			10'd528: USel4 = 4'b0100;
			10'd529: USel4 = 4'b0100;
			10'd530: USel4 = 4'b1000;
			10'd531: USel4 = 4'b1000;
			10'd532: USel4 = 4'b1000;
			10'd533: USel4 = 4'b1000;
			10'd534: USel4 = 4'b1000;
			10'd535: USel4 = 4'b1000;
			10'd536: USel4 = 4'b1000;
			10'd537: USel4 = 4'b1000;
			10'd538: USel4 = 4'b1000;
			10'd539: USel4 = 4'b1000;
			10'd540: USel4 = 4'b1000;
			10'd541: USel4 = 4'b1000;
			10'd542: USel4 = 4'b1000;
			10'd543: USel4 = 4'b1000;
			10'd544: USel4 = 4'b1000;
			10'd545: USel4 = 4'b1000;
			10'd546: USel4 = 4'b1000;
			10'd547: USel4 = 4'b1000;
			10'd548: USel4 = 4'b1000;
			10'd549: USel4 = 4'b1000;
			10'd550: USel4 = 4'b1000;
			10'd551: USel4 = 4'b1000;
			10'd552: USel4 = 4'b1000;
			10'd553: USel4 = 4'b1000;
			10'd554: USel4 = 4'b1000;
			10'd555: USel4 = 4'b1000;
			10'd556: USel4 = 4'b1000;
			10'd557: USel4 = 4'b1000;
			10'd558: USel4 = 4'b1000;
			10'd559: USel4 = 4'b1000;
			10'd560: USel4 = 4'b1000;
			10'd561: USel4 = 4'b1000;
			10'd562: USel4 = 4'b1000;
			10'd563: USel4 = 4'b1000;
			10'd564: USel4 = 4'b1000;
			10'd565: USel4 = 4'b1000;
			10'd566: USel4 = 4'b1000;
			10'd567: USel4 = 4'b1000;
			10'd568: USel4 = 4'b1000;
			10'd569: USel4 = 4'b1000;
			10'd570: USel4 = 4'b1000;
			10'd571: USel4 = 4'b1000;
			10'd572: USel4 = 4'b1000;
			10'd573: USel4 = 4'b1000;
			10'd574: USel4 = 4'b1000;
			10'd575: USel4 = 4'b1000;
			10'd576: USel4 = 4'b0001;
			10'd577: USel4 = 4'b0001;
			10'd578: USel4 = 4'b0001;
			10'd579: USel4 = 4'b0001;
			10'd580: USel4 = 4'b0001;
			10'd581: USel4 = 4'b0001;
			10'd582: USel4 = 4'b0001;
			10'd583: USel4 = 4'b0001;
			10'd584: USel4 = 4'b0001;
			10'd585: USel4 = 4'b0001;
			10'd586: USel4 = 4'b0001;
			10'd587: USel4 = 4'b0001;
			10'd588: USel4 = 4'b0001;
			10'd589: USel4 = 4'b0001;
			10'd590: USel4 = 4'b0001;
			10'd591: USel4 = 4'b0001;
			10'd592: USel4 = 4'b0001;
			10'd593: USel4 = 4'b0001;
			10'd594: USel4 = 4'b0001;
			10'd595: USel4 = 4'b0001;
			10'd596: USel4 = 4'b0001;
			10'd597: USel4 = 4'b0001;
			10'd598: USel4 = 4'b0001;
			10'd599: USel4 = 4'b0001;
			10'd600: USel4 = 4'b0001;
			10'd601: USel4 = 4'b0001;
			10'd602: USel4 = 4'b0001;
			10'd603: USel4 = 4'b0001;
			10'd604: USel4 = 4'b0001;
			10'd605: USel4 = 4'b0001;
			10'd606: USel4 = 4'b0001;
			10'd607: USel4 = 4'b0001;
			10'd608: USel4 = 4'b0001;
			10'd609: USel4 = 4'b0001;
			10'd610: USel4 = 4'b0001;
			10'd611: USel4 = 4'b0001;
			10'd612: USel4 = 4'b0001;
			10'd613: USel4 = 4'b0001;
			10'd614: USel4 = 4'b0001;
			10'd615: USel4 = 4'b0001;
			10'd616: USel4 = 4'b0001;
			10'd617: USel4 = 4'b0001;
			10'd618: USel4 = 4'b0001;
			10'd619: USel4 = 4'b0001;
			10'd620: USel4 = 4'b0001;
			10'd621: USel4 = 4'b0001;
			10'd622: USel4 = 4'b0010;
			10'd623: USel4 = 4'b0010;
			10'd624: USel4 = 4'b0010;
			10'd625: USel4 = 4'b0010;
			10'd626: USel4 = 4'b0010;
			10'd627: USel4 = 4'b0010;
			10'd628: USel4 = 4'b0010;
			10'd629: USel4 = 4'b0010;
			10'd630: USel4 = 4'b0010;
			10'd631: USel4 = 4'b0010;
			10'd632: USel4 = 4'b0010;
			10'd633: USel4 = 4'b0010;
			10'd634: USel4 = 4'b0000;
			10'd635: USel4 = 4'b0000;
			10'd636: USel4 = 4'b0000;
			10'd637: USel4 = 4'b0000;
			10'd638: USel4 = 4'b0000;
			10'd639: USel4 = 4'b0000;
			10'd640: USel4 = 4'b0000;
			10'd641: USel4 = 4'b0000;
			10'd642: USel4 = 4'b0000;
			10'd643: USel4 = 4'b0000;
			10'd644: USel4 = 4'b0000;
			10'd645: USel4 = 4'b0000;
			10'd646: USel4 = 4'b0100;
			10'd647: USel4 = 4'b0100;
			10'd648: USel4 = 4'b0100;
			10'd649: USel4 = 4'b0100;
			10'd650: USel4 = 4'b0100;
			10'd651: USel4 = 4'b0100;
			10'd652: USel4 = 4'b0100;
			10'd653: USel4 = 4'b0100;
			10'd654: USel4 = 4'b0100;
			10'd655: USel4 = 4'b0100;
			10'd656: USel4 = 4'b0100;
			10'd657: USel4 = 4'b0100;
			10'd658: USel4 = 4'b0100;
			10'd659: USel4 = 4'b0100;
			10'd660: USel4 = 4'b1000;
			10'd661: USel4 = 4'b1000;
			10'd662: USel4 = 4'b1000;
			10'd663: USel4 = 4'b1000;
			10'd664: USel4 = 4'b1000;
			10'd665: USel4 = 4'b1000;
			10'd666: USel4 = 4'b1000;
			10'd667: USel4 = 4'b1000;
			10'd668: USel4 = 4'b1000;
			10'd669: USel4 = 4'b1000;
			10'd670: USel4 = 4'b1000;
			10'd671: USel4 = 4'b1000;
			10'd672: USel4 = 4'b1000;
			10'd673: USel4 = 4'b1000;
			10'd674: USel4 = 4'b1000;
			10'd675: USel4 = 4'b1000;
			10'd676: USel4 = 4'b1000;
			10'd677: USel4 = 4'b1000;
			10'd678: USel4 = 4'b1000;
			10'd679: USel4 = 4'b1000;
			10'd680: USel4 = 4'b1000;
			10'd681: USel4 = 4'b1000;
			10'd682: USel4 = 4'b1000;
			10'd683: USel4 = 4'b1000;
			10'd684: USel4 = 4'b1000;
			10'd685: USel4 = 4'b1000;
			10'd686: USel4 = 4'b1000;
			10'd687: USel4 = 4'b1000;
			10'd688: USel4 = 4'b1000;
			10'd689: USel4 = 4'b1000;
			10'd690: USel4 = 4'b1000;
			10'd691: USel4 = 4'b1000;
			10'd692: USel4 = 4'b1000;
			10'd693: USel4 = 4'b1000;
			10'd694: USel4 = 4'b1000;
			10'd695: USel4 = 4'b1000;
			10'd696: USel4 = 4'b1000;
			10'd697: USel4 = 4'b1000;
			10'd698: USel4 = 4'b1000;
			10'd699: USel4 = 4'b1000;
			10'd700: USel4 = 4'b1000;
			10'd701: USel4 = 4'b1000;
			10'd702: USel4 = 4'b1000;
			10'd703: USel4 = 4'b1000;
			10'd704: USel4 = 4'b0001;
			10'd705: USel4 = 4'b0001;
			10'd706: USel4 = 4'b0001;
			10'd707: USel4 = 4'b0001;
			10'd708: USel4 = 4'b0001;
			10'd709: USel4 = 4'b0001;
			10'd710: USel4 = 4'b0001;
			10'd711: USel4 = 4'b0001;
			10'd712: USel4 = 4'b0001;
			10'd713: USel4 = 4'b0001;
			10'd714: USel4 = 4'b0001;
			10'd715: USel4 = 4'b0001;
			10'd716: USel4 = 4'b0001;
			10'd717: USel4 = 4'b0001;
			10'd718: USel4 = 4'b0001;
			10'd719: USel4 = 4'b0001;
			10'd720: USel4 = 4'b0001;
			10'd721: USel4 = 4'b0001;
			10'd722: USel4 = 4'b0001;
			10'd723: USel4 = 4'b0001;
			10'd724: USel4 = 4'b0001;
			10'd725: USel4 = 4'b0001;
			10'd726: USel4 = 4'b0001;
			10'd727: USel4 = 4'b0001;
			10'd728: USel4 = 4'b0001;
			10'd729: USel4 = 4'b0001;
			10'd730: USel4 = 4'b0001;
			10'd731: USel4 = 4'b0001;
			10'd732: USel4 = 4'b0001;
			10'd733: USel4 = 4'b0001;
			10'd734: USel4 = 4'b0001;
			10'd735: USel4 = 4'b0001;
			10'd736: USel4 = 4'b0001;
			10'd737: USel4 = 4'b0001;
			10'd738: USel4 = 4'b0001;
			10'd739: USel4 = 4'b0001;
			10'd740: USel4 = 4'b0001;
			10'd741: USel4 = 4'b0001;
			10'd742: USel4 = 4'b0001;
			10'd743: USel4 = 4'b0001;
			10'd744: USel4 = 4'b0001;
			10'd745: USel4 = 4'b0001;
			10'd746: USel4 = 4'b0001;
			10'd747: USel4 = 4'b0001;
			10'd748: USel4 = 4'b0010;
			10'd749: USel4 = 4'b0010;
			10'd750: USel4 = 4'b0010;
			10'd751: USel4 = 4'b0010;
			10'd752: USel4 = 4'b0010;
			10'd753: USel4 = 4'b0010;
			10'd754: USel4 = 4'b0010;
			10'd755: USel4 = 4'b0010;
			10'd756: USel4 = 4'b0010;
			10'd757: USel4 = 4'b0010;
			10'd758: USel4 = 4'b0010;
			10'd759: USel4 = 4'b0010;
			10'd760: USel4 = 4'b0000;
			10'd761: USel4 = 4'b0000;
			10'd762: USel4 = 4'b0000;
			10'd763: USel4 = 4'b0000;
			10'd764: USel4 = 4'b0000;
			10'd765: USel4 = 4'b0000;
			10'd766: USel4 = 4'b0000;
			10'd767: USel4 = 4'b0000;
			10'd768: USel4 = 4'b0000;
			10'd769: USel4 = 4'b0000;
			10'd770: USel4 = 4'b0000;
			10'd771: USel4 = 4'b0000;
			10'd772: USel4 = 4'b0000;
			10'd773: USel4 = 4'b0000;
			10'd774: USel4 = 4'b0000;
			10'd775: USel4 = 4'b0000;
			10'd776: USel4 = 4'b0100;
			10'd777: USel4 = 4'b0100;
			10'd778: USel4 = 4'b0100;
			10'd779: USel4 = 4'b0100;
			10'd780: USel4 = 4'b0100;
			10'd781: USel4 = 4'b0100;
			10'd782: USel4 = 4'b0100;
			10'd783: USel4 = 4'b0100;
			10'd784: USel4 = 4'b0100;
			10'd785: USel4 = 4'b0100;
			10'd786: USel4 = 4'b0100;
			10'd787: USel4 = 4'b0100;
			10'd788: USel4 = 4'b1000;
			10'd789: USel4 = 4'b1000;
			10'd790: USel4 = 4'b1000;
			10'd791: USel4 = 4'b1000;
			10'd792: USel4 = 4'b1000;
			10'd793: USel4 = 4'b1000;
			10'd794: USel4 = 4'b1000;
			10'd795: USel4 = 4'b1000;
			10'd796: USel4 = 4'b1000;
			10'd797: USel4 = 4'b1000;
			10'd798: USel4 = 4'b1000;
			10'd799: USel4 = 4'b1000;
			10'd800: USel4 = 4'b1000;
			10'd801: USel4 = 4'b1000;
			10'd802: USel4 = 4'b1000;
			10'd803: USel4 = 4'b1000;
			10'd804: USel4 = 4'b1000;
			10'd805: USel4 = 4'b1000;
			10'd806: USel4 = 4'b1000;
			10'd807: USel4 = 4'b1000;
			10'd808: USel4 = 4'b1000;
			10'd809: USel4 = 4'b1000;
			10'd810: USel4 = 4'b1000;
			10'd811: USel4 = 4'b1000;
			10'd812: USel4 = 4'b1000;
			10'd813: USel4 = 4'b1000;
			10'd814: USel4 = 4'b1000;
			10'd815: USel4 = 4'b1000;
			10'd816: USel4 = 4'b1000;
			10'd817: USel4 = 4'b1000;
			10'd818: USel4 = 4'b1000;
			10'd819: USel4 = 4'b1000;
			10'd820: USel4 = 4'b1000;
			10'd821: USel4 = 4'b1000;
			10'd822: USel4 = 4'b1000;
			10'd823: USel4 = 4'b1000;
			10'd824: USel4 = 4'b1000;
			10'd825: USel4 = 4'b1000;
			10'd826: USel4 = 4'b1000;
			10'd827: USel4 = 4'b1000;
			10'd828: USel4 = 4'b1000;
			10'd829: USel4 = 4'b1000;
			10'd830: USel4 = 4'b1000;
			10'd831: USel4 = 4'b1000;
			10'd832: USel4 = 4'b0001;
			10'd833: USel4 = 4'b0001;
			10'd834: USel4 = 4'b0001;
			10'd835: USel4 = 4'b0001;
			10'd836: USel4 = 4'b0001;
			10'd837: USel4 = 4'b0001;
			10'd838: USel4 = 4'b0001;
			10'd839: USel4 = 4'b0001;
			10'd840: USel4 = 4'b0001;
			10'd841: USel4 = 4'b0001;
			10'd842: USel4 = 4'b0001;
			10'd843: USel4 = 4'b0001;
			10'd844: USel4 = 4'b0001;
			10'd845: USel4 = 4'b0001;
			10'd846: USel4 = 4'b0001;
			10'd847: USel4 = 4'b0001;
			10'd848: USel4 = 4'b0001;
			10'd849: USel4 = 4'b0001;
			10'd850: USel4 = 4'b0001;
			10'd851: USel4 = 4'b0001;
			10'd852: USel4 = 4'b0001;
			10'd853: USel4 = 4'b0001;
			10'd854: USel4 = 4'b0001;
			10'd855: USel4 = 4'b0001;
			10'd856: USel4 = 4'b0001;
			10'd857: USel4 = 4'b0001;
			10'd858: USel4 = 4'b0001;
			10'd859: USel4 = 4'b0001;
			10'd860: USel4 = 4'b0001;
			10'd861: USel4 = 4'b0001;
			10'd862: USel4 = 4'b0001;
			10'd863: USel4 = 4'b0001;
			10'd864: USel4 = 4'b0001;
			10'd865: USel4 = 4'b0001;
			10'd866: USel4 = 4'b0001;
			10'd867: USel4 = 4'b0001;
			10'd868: USel4 = 4'b0001;
			10'd869: USel4 = 4'b0001;
			10'd870: USel4 = 4'b0001;
			10'd871: USel4 = 4'b0001;
			10'd872: USel4 = 4'b0001;
			10'd873: USel4 = 4'b0001;
			10'd874: USel4 = 4'b0010;
			10'd875: USel4 = 4'b0010;
			10'd876: USel4 = 4'b0010;
			10'd877: USel4 = 4'b0010;
			10'd878: USel4 = 4'b0010;
			10'd879: USel4 = 4'b0010;
			10'd880: USel4 = 4'b0010;
			10'd881: USel4 = 4'b0010;
			10'd882: USel4 = 4'b0010;
			10'd883: USel4 = 4'b0010;
			10'd884: USel4 = 4'b0010;
			10'd885: USel4 = 4'b0010;
			10'd886: USel4 = 4'b0010;
			10'd887: USel4 = 4'b0010;
			10'd888: USel4 = 4'b0000;
			10'd889: USel4 = 4'b0000;
			10'd890: USel4 = 4'b0000;
			10'd891: USel4 = 4'b0000;
			10'd892: USel4 = 4'b0000;
			10'd893: USel4 = 4'b0000;
			10'd894: USel4 = 4'b0000;
			10'd895: USel4 = 4'b0000;
			10'd896: USel4 = 4'b0000;
			10'd897: USel4 = 4'b0000;
			10'd898: USel4 = 4'b0000;
			10'd899: USel4 = 4'b0000;
			10'd900: USel4 = 4'b0000;
			10'd901: USel4 = 4'b0000;
			10'd902: USel4 = 4'b0000;
			10'd903: USel4 = 4'b0000;
			10'd904: USel4 = 4'b0100;
			10'd905: USel4 = 4'b0100;
			10'd906: USel4 = 4'b0100;
			10'd907: USel4 = 4'b0100;
			10'd908: USel4 = 4'b0100;
			10'd909: USel4 = 4'b0100;
			10'd910: USel4 = 4'b0100;
			10'd911: USel4 = 4'b0100;
			10'd912: USel4 = 4'b0100;
			10'd913: USel4 = 4'b0100;
			10'd914: USel4 = 4'b0100;
			10'd915: USel4 = 4'b0100;
			10'd916: USel4 = 4'b0100;
			10'd917: USel4 = 4'b0100;
			10'd918: USel4 = 4'b0100;
			10'd919: USel4 = 4'b0100;
			10'd920: USel4 = 4'b1000;
			10'd921: USel4 = 4'b1000;
			10'd922: USel4 = 4'b1000;
			10'd923: USel4 = 4'b1000;
			10'd924: USel4 = 4'b1000;
			10'd925: USel4 = 4'b1000;
			10'd926: USel4 = 4'b1000;
			10'd927: USel4 = 4'b1000;
			10'd928: USel4 = 4'b1000;
			10'd929: USel4 = 4'b1000;
			10'd930: USel4 = 4'b1000;
			10'd931: USel4 = 4'b1000;
			10'd932: USel4 = 4'b1000;
			10'd933: USel4 = 4'b1000;
			10'd934: USel4 = 4'b1000;
			10'd935: USel4 = 4'b1000;
			10'd936: USel4 = 4'b1000;
			10'd937: USel4 = 4'b1000;
			10'd938: USel4 = 4'b1000;
			10'd939: USel4 = 4'b1000;
			10'd940: USel4 = 4'b1000;
			10'd941: USel4 = 4'b1000;
			10'd942: USel4 = 4'b1000;
			10'd943: USel4 = 4'b1000;
			10'd944: USel4 = 4'b1000;
			10'd945: USel4 = 4'b1000;
			10'd946: USel4 = 4'b1000;
			10'd947: USel4 = 4'b1000;
			10'd948: USel4 = 4'b1000;
			10'd949: USel4 = 4'b1000;
			10'd950: USel4 = 4'b1000;
			10'd951: USel4 = 4'b1000;
			10'd952: USel4 = 4'b1000;
			10'd953: USel4 = 4'b1000;
			10'd954: USel4 = 4'b1000;
			10'd955: USel4 = 4'b1000;
			10'd956: USel4 = 4'b1000;
			10'd957: USel4 = 4'b1000;
			10'd958: USel4 = 4'b1000;
			10'd959: USel4 = 4'b1000;
			10'd960: USel4 = 4'b0001;
			10'd961: USel4 = 4'b0001;
			10'd962: USel4 = 4'b0001;
			10'd963: USel4 = 4'b0001;
			10'd964: USel4 = 4'b0001;
			10'd965: USel4 = 4'b0001;
			10'd966: USel4 = 4'b0001;
			10'd967: USel4 = 4'b0001;
			10'd968: USel4 = 4'b0001;
			10'd969: USel4 = 4'b0001;
			10'd970: USel4 = 4'b0001;
			10'd971: USel4 = 4'b0001;
			10'd972: USel4 = 4'b0001;
			10'd973: USel4 = 4'b0001;
			10'd974: USel4 = 4'b0001;
			10'd975: USel4 = 4'b0001;
			10'd976: USel4 = 4'b0001;
			10'd977: USel4 = 4'b0001;
			10'd978: USel4 = 4'b0001;
			10'd979: USel4 = 4'b0001;
			10'd980: USel4 = 4'b0001;
			10'd981: USel4 = 4'b0001;
			10'd982: USel4 = 4'b0001;
			10'd983: USel4 = 4'b0001;
			10'd984: USel4 = 4'b0001;
			10'd985: USel4 = 4'b0001;
			10'd986: USel4 = 4'b0001;
			10'd987: USel4 = 4'b0001;
			10'd988: USel4 = 4'b0001;
			10'd989: USel4 = 4'b0001;
			10'd990: USel4 = 4'b0001;
			10'd991: USel4 = 4'b0001;
			10'd992: USel4 = 4'b0001;
			10'd993: USel4 = 4'b0001;
			10'd994: USel4 = 4'b0001;
			10'd995: USel4 = 4'b0001;
			10'd996: USel4 = 4'b0001;
			10'd997: USel4 = 4'b0001;
			10'd998: USel4 = 4'b0001;
			10'd999: USel4 = 4'b0001;
			10'd1000: USel4 = 4'b0001;
			10'd1001: USel4 = 4'b0001;
			10'd1002: USel4 = 4'b0010;
			10'd1003: USel4 = 4'b0010;
			10'd1004: USel4 = 4'b0010;
			10'd1005: USel4 = 4'b0010;
			10'd1006: USel4 = 4'b0010;
			10'd1007: USel4 = 4'b0010;
			10'd1008: USel4 = 4'b0010;
			10'd1009: USel4 = 4'b0010;
			10'd1010: USel4 = 4'b0010;
			10'd1011: USel4 = 4'b0010;
			10'd1012: USel4 = 4'b0010;
			10'd1013: USel4 = 4'b0010;
			10'd1014: USel4 = 4'b0010;
			10'd1015: USel4 = 4'b0010;
			10'd1016: USel4 = 4'b0000;
			10'd1017: USel4 = 4'b0000;
			10'd1018: USel4 = 4'b0000;
			10'd1019: USel4 = 4'b0000;
			10'd1020: USel4 = 4'b0000;
			10'd1021: USel4 = 4'b0000;
			10'd1022: USel4 = 4'b0000;
			10'd1023: USel4 = 4'b0000;
		endcase
	end
	always @(*) begin
		if (_sv2v_0)
			;
		if (Sqrt) begin
			if (j1)
				A = 3'b101;
			else if (Smsbs[4] == 1)
				A = 3'b111;
			else
				A = Smsbs[2:0];
		end
		else
			A = Dmsbs;
	end
	assign udigit = (Sqrt & j0 ? 4'b0100 : USel4);
	initial _sv2v_0 = 0;
endmodule
module fma (
	Xs,
	Ys,
	Zs,
	Xe,
	Ye,
	Ze,
	Xm,
	Ym,
	Zm,
	XZero,
	YZero,
	ZZero,
	OpCtrl,
	ASticky,
	Sm,
	InvA,
	As,
	Ps,
	Ss,
	Se,
	SCnt
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire Xs;
	input wire Ys;
	input wire Zs;
	input wire [$signed(P[837-:32]) - 1:0] Xe;
	input wire [$signed(P[837-:32]) - 1:0] Ye;
	input wire [$signed(P[837-:32]) - 1:0] Ze;
	input wire [$signed(P[805-:32]):0] Xm;
	input wire [$signed(P[805-:32]):0] Ym;
	input wire [$signed(P[805-:32]):0] Zm;
	input wire XZero;
	input wire YZero;
	input wire ZZero;
	input wire [2:0] OpCtrl;
	output wire ASticky;
	output wire [$signed(P[255-:32]) - 1:0] Sm;
	output wire InvA;
	output wire As;
	output wire Ps;
	output wire Ss;
	output wire [$signed(P[837-:32]) + 1:0] Se;
	output wire [$clog2($signed(P[255-:32]) + 1) - 1:0] SCnt;
	wire [(2 * $signed(P[805-:32])) + 1:0] Pm;
	wire [$signed(P[255-:32]) - 1:0] Am;
	wire [$signed(P[255-:32]) - 1:0] AmInv;
	wire [(2 * $signed(P[805-:32])) + 1:0] PmKilled;
	wire KillProd;
	wire [$signed(P[837-:32]) + 1:0] Pe;
	fmaexpadd #(.P(P)) expadd(
		.Xe(Xe),
		.Ye(Ye),
		.XZero(XZero),
		.YZero(YZero),
		.Pe(Pe)
	);
	fmamult #(.P(P)) mult(
		.Xm(Xm),
		.Ym(Ym),
		.Pm(Pm)
	);
	fmasign sign(
		.OpCtrl(OpCtrl),
		.Xs(Xs),
		.Ys(Ys),
		.Zs(Zs),
		.Ps(Ps),
		.As(As),
		.InvA(InvA)
	);
	fmaalign #(.P(P)) align(
		.Ze(Ze),
		.Zm(Zm),
		.XZero(XZero),
		.YZero(YZero),
		.ZZero(ZZero),
		.Xe(Xe),
		.Ye(Ye),
		.Am(Am),
		.ASticky(ASticky),
		.KillProd(KillProd)
	);
	fmaadd #(.P(P)) add(
		.Am(Am),
		.Pm(Pm),
		.Ze(Ze),
		.Pe(Pe),
		.Ps(Ps),
		.KillProd(KillProd),
		.ASticky(ASticky),
		.AmInv(AmInv),
		.PmKilled(PmKilled),
		.InvA(InvA),
		.Sm(Sm),
		.Se(Se),
		.Ss(Ss)
	);
	fmalza #(
		.WIDTH($signed(P[255-:32])),
		.NF($signed(P[805-:32]))
	) lza(
		.A(AmInv),
		.Pm(PmKilled),
		.Cin(InvA & (~ASticky | KillProd)),
		.sub(InvA),
		.SCnt(SCnt)
	);
endmodule
module fmaadd (
	Am,
	Ze,
	Ps,
	Pe,
	Pm,
	InvA,
	KillProd,
	ASticky,
	AmInv,
	PmKilled,
	Ss,
	Se,
	Sm
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [(3 * $signed(P[805-:32])) + 5:0] Am;
	input wire [$signed(P[837-:32]) - 1:0] Ze;
	input wire Ps;
	input wire [$signed(P[837-:32]) + 1:0] Pe;
	input wire [(2 * $signed(P[805-:32])) + 1:0] Pm;
	input wire InvA;
	input wire KillProd;
	input wire ASticky;
	output wire [(3 * $signed(P[805-:32])) + 5:0] AmInv;
	output wire [(2 * $signed(P[805-:32])) + 1:0] PmKilled;
	output wire Ss;
	output wire [$signed(P[837-:32]) + 1:0] Se;
	output wire [(3 * $signed(P[805-:32])) + 5:0] Sm;
	wire [(3 * $signed(P[805-:32])) + 5:0] PreSum;
	wire [(3 * $signed(P[805-:32])) + 5:0] NegPreSum;
	wire NegSum;
	assign AmInv = (InvA ? ~Am : Am);
	assign PmKilled = (KillProd ? 0 : Pm);
	assign {NegSum, PreSum} = ({{$signed(P[805-:32]) + 3 {1'b0}}, PmKilled, 2'b00} + {InvA, AmInv}) + {{(3 * $signed(P[805-:32])) + 5 {1'b0}}, (~ASticky | KillProd) & InvA};
	function automatic signed [(((3 * $signed(P[805-:32])) + 2) >= 0 ? (3 * $signed(P[805-:32])) + 3 : 1 - ((3 * $signed(P[805-:32])) + 2)) - 1:0] sv2v_cast_B52D7_signed;
		input reg signed [(((3 * $signed(P[805-:32])) + 2) >= 0 ? (3 * $signed(P[805-:32])) + 3 : 1 - ((3 * $signed(P[805-:32])) + 2)) - 1:0] inp;
		sv2v_cast_B52D7_signed = inp;
	endfunction
	assign NegPreSum = (Am + {{$signed(P[805-:32]) + 2 {1'b1}}, ~PmKilled, 2'b00}) + {sv2v_cast_B52D7_signed(0), ~ASticky | ~KillProd, 2'b00};
	assign Sm = (NegSum ? NegPreSum : PreSum);
	assign Ss = NegSum ^ Ps;
	assign Se = (KillProd ? {2'b00, Ze} : Pe);
endmodule
module fmaalign (
	Xe,
	Ye,
	Ze,
	Zm,
	XZero,
	YZero,
	ZZero,
	Am,
	ASticky,
	KillProd
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[837-:32]) - 1:0] Xe;
	input wire [$signed(P[837-:32]) - 1:0] Ye;
	input wire [$signed(P[837-:32]) - 1:0] Ze;
	input wire [$signed(P[805-:32]):0] Zm;
	input wire XZero;
	input wire YZero;
	input wire ZZero;
	output wire [$signed(P[255-:32]) - 1:0] Am;
	output reg ASticky;
	output wire KillProd;
	wire [$signed(P[837-:32]) + 1:0] ACnt;
	reg [($signed(P[255-:32]) + $signed(P[805-:32])) - 1:0] ZmShifted;
	wire [($signed(P[255-:32]) + $signed(P[805-:32])) - 1:0] ZmPreshifted;
	wire KillZ;
	function automatic signed [$signed(P[837-:32]) - 1:0] sv2v_cast_AF3D4_signed;
		input reg signed [$signed(P[837-:32]) - 1:0] inp;
		sv2v_cast_AF3D4_signed = inp;
	endfunction
	function automatic signed [(($signed(P[837-:32]) + 1) >= 0 ? $signed(P[837-:32]) + 2 : 1 - ($signed(P[837-:32]) + 1)) - 1:0] sv2v_cast_A1EFF_signed;
		input reg signed [(($signed(P[837-:32]) + 1) >= 0 ? $signed(P[837-:32]) + 2 : 1 - ($signed(P[837-:32]) + 1)) - 1:0] inp;
		sv2v_cast_A1EFF_signed = inp;
	endfunction
	assign ACnt = ((({2'b00, Xe} + {2'b00, Ye}) - {2'b00, sv2v_cast_AF3D4_signed($signed(P[771-:32]))}) + sv2v_cast_A1EFF_signed($signed(P[805-:32]) + 3)) - {2'b00, Ze};
	function automatic signed [(($signed(P[255-:32]) - 2) >= 0 ? $signed(P[255-:32]) - 1 : 3 - $signed(P[255-:32])) - 1:0] sv2v_cast_1AFFE_signed;
		input reg signed [(($signed(P[255-:32]) - 2) >= 0 ? $signed(P[255-:32]) - 1 : 3 - $signed(P[255-:32])) - 1:0] inp;
		sv2v_cast_1AFFE_signed = inp;
	endfunction
	assign ZmPreshifted = {Zm, sv2v_cast_1AFFE_signed(0)};
	assign KillProd = ((ACnt[$signed(P[837-:32]) + 1] & ~ZZero) | XZero) | YZero;
	assign KillZ = $signed(ACnt) > $signed((sv2v_cast_A1EFF_signed(3) * sv2v_cast_A1EFF_signed($signed(P[805-:32]))) + sv2v_cast_A1EFF_signed(5));
	function automatic signed [(($signed(P[805-:32]) + 2) >= 0 ? $signed(P[805-:32]) + 3 : 1 - ($signed(P[805-:32]) + 2)) - 1:0] sv2v_cast_BC2DD_signed;
		input reg signed [(($signed(P[805-:32]) + 2) >= 0 ? $signed(P[805-:32]) + 3 : 1 - ($signed(P[805-:32]) + 2)) - 1:0] inp;
		sv2v_cast_BC2DD_signed = inp;
	endfunction
	function automatic signed [(((2 * $signed(P[805-:32])) + 1) >= 0 ? (2 * $signed(P[805-:32])) + 2 : 1 - ((2 * $signed(P[805-:32])) + 1)) - 1:0] sv2v_cast_C99B7_signed;
		input reg signed [(((2 * $signed(P[805-:32])) + 1) >= 0 ? (2 * $signed(P[805-:32])) + 2 : 1 - ((2 * $signed(P[805-:32])) + 1)) - 1:0] inp;
		sv2v_cast_C99B7_signed = inp;
	endfunction
	always @(*) begin
		if (_sv2v_0)
			;
		if (KillProd) begin
			ZmShifted = {sv2v_cast_BC2DD_signed(0), Zm, sv2v_cast_C99B7_signed(0)};
			ASticky = ~(XZero | YZero);
		end
		else if (KillZ) begin
			ZmShifted = 1'sb0;
			ASticky = ~ZZero;
		end
		else begin
			ZmShifted = ZmPreshifted >> ACnt;
			ASticky = |ZmShifted[$signed(P[805-:32]) - 1:0];
		end
	end
	assign Am = ZmShifted[($signed(P[255-:32]) + $signed(P[805-:32])) - 1:$signed(P[805-:32])];
	initial _sv2v_0 = 0;
endmodule
module fmaexpadd (
	Xe,
	Ye,
	XZero,
	YZero,
	Pe
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[837-:32]) - 1:0] Xe;
	input wire [$signed(P[837-:32]) - 1:0] Ye;
	input wire XZero;
	input wire YZero;
	output wire [$signed(P[837-:32]) + 1:0] Pe;
	wire PZero;
	assign PZero = XZero | YZero;
	function automatic signed [$signed(P[837-:32]) - 1:0] sv2v_cast_AF3D4_signed;
		input reg signed [$signed(P[837-:32]) - 1:0] inp;
		sv2v_cast_AF3D4_signed = inp;
	endfunction
	assign Pe = (PZero ? {(($signed(P[837-:32]) + 1) >= 0 ? $signed(P[837-:32]) + 2 : 1 - ($signed(P[837-:32]) + 1)) {1'sb0}} : ({2'b00, Xe} + {2'b00, Ye}) - {2'b00, sv2v_cast_AF3D4_signed($signed(P[771-:32]))});
endmodule
module fmalza (
	A,
	Pm,
	Cin,
	sub,
	SCnt
);
	parameter WIDTH = 0;
	parameter NF = 0;
	input wire [WIDTH - 1:0] A;
	input wire [(2 * NF) + 1:0] Pm;
	input wire Cin;
	input wire sub;
	output wire [$clog2(WIDTH + 1) - 1:0] SCnt;
	wire [WIDTH:0] F;
	wire [WIDTH - 1:0] B;
	wire [WIDTH - 1:0] P;
	wire [WIDTH - 1:0] G;
	wire [WIDTH - 1:0] K;
	wire [WIDTH - 1:0] Pp1;
	wire [WIDTH - 1:0] Gm1;
	wire [WIDTH - 1:0] Km1;
	assign B = {{NF + 2 {1'b0}}, Pm, 2'b00};
	assign P = A ^ B;
	assign G = A & B;
	assign K = ~A & ~B;
	assign Pp1 = {sub, P[WIDTH - 1:1]};
	assign Gm1 = {G[WIDTH - 2:0], Cin};
	assign Km1 = {K[WIDTH - 2:0], ~Cin};
	assign F[WIDTH] = ~sub & P[WIDTH - 1];
	assign F[WIDTH - 1:0] = (Pp1 & ((G & ~Km1) | (K & ~Gm1))) | (~Pp1 & ((K & ~Km1) | (G & ~Gm1)));
	lzc #(.WIDTH(WIDTH + 1)) lzc(
		.num(F),
		.ZeroCnt(SCnt)
	);
endmodule
module fmamult (
	Xm,
	Ym,
	Pm
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[805-:32]):0] Xm;
	input wire [$signed(P[805-:32]):0] Ym;
	output wire [(2 * $signed(P[805-:32])) + 1:0] Pm;
	assign Pm = Xm * Ym;
endmodule
module fmasign (
	OpCtrl,
	Xs,
	Ys,
	Zs,
	Ps,
	As,
	InvA
);
	input wire [2:0] OpCtrl;
	input wire Xs;
	input wire Ys;
	input wire Zs;
	output wire Ps;
	output wire As;
	output wire InvA;
	assign Ps = (Xs ^ Ys) ^ (OpCtrl[1] & ~OpCtrl[2]);
	assign As = Zs ^ OpCtrl[0];
	assign InvA = As ^ Ps;
endmodule
module cvtshiftcalc (
	XZero,
	ToInt,
	IntToFp,
	OutFmt,
	CvtCe,
	Xm,
	CvtLzcIn,
	CvtResSubnormUf,
	CvtResUf,
	CvtShiftIn
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire XZero;
	input wire ToInt;
	input wire IntToFp;
	input wire [$signed(P[707-:32]) - 1:0] OutFmt;
	input wire [$signed(P[837-:32]):0] CvtCe;
	input wire [$signed(P[805-:32]):0] Xm;
	input wire [$signed(P[415-:32]) - 1:0] CvtLzcIn;
	input wire CvtResSubnormUf;
	output wire CvtResUf;
	output reg [$signed(P[415-:32]) + $signed(P[805-:32]):0] CvtShiftIn;
	reg [$clog2($signed(P[805-:32])):0] ResNegNF;
	always @(*) begin
		if (_sv2v_0)
			;
		if (ToInt)
			CvtShiftIn = {{$signed(P[4216-:32]) {1'b0}}, Xm[$signed(P[805-:32])] & ~CvtCe[$signed(P[837-:32])], Xm[$signed(P[805-:32]) - 1] | (CvtCe[$signed(P[837-:32])] & Xm[$signed(P[805-:32])]), Xm[$signed(P[805-:32]) - 2:0], {$signed(P[415-:32]) - $signed(P[4216-:32]) {1'b0}}};
		else if (CvtResSubnormUf)
			CvtShiftIn = {{$signed(P[805-:32]) - 1 {1'b0}}, Xm, {($signed(P[415-:32]) - $signed(P[805-:32])) + 1 {1'b0}}};
		else
			CvtShiftIn = {CvtLzcIn, {$signed(P[805-:32]) + 1 {1'b0}}};
	end
	function automatic signed [(($clog2($signed(P[805-:32])) + 0) >= 0 ? $clog2($signed(P[805-:32])) + 1 : 1 - ($clog2($signed(P[805-:32])) + 0)) - 1:0] sv2v_cast_D43F7_signed;
		input reg signed [(($clog2($signed(P[805-:32])) + 0) >= 0 ? $clog2($signed(P[805-:32])) + 1 : 1 - ($clog2($signed(P[805-:32])) + 0)) - 1:0] inp;
		sv2v_cast_D43F7_signed = inp;
	endfunction
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk1
			wire [($clog2($signed(P[805-:32])) >= 0 ? $clog2($signed(P[805-:32])) + 1 : 1 - $clog2($signed(P[805-:32]))):1] sv2v_tmp_9FF21;
			assign sv2v_tmp_9FF21 = -sv2v_cast_D43F7_signed($signed(P[805-:32]));
			always @(*) ResNegNF = sv2v_tmp_9FF21;
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk1
			wire [($clog2($signed(P[805-:32])) >= 0 ? $clog2($signed(P[805-:32])) + 1 : 1 - $clog2($signed(P[805-:32]))):1] sv2v_tmp_DB608;
			assign sv2v_tmp_DB608 = (OutFmt ? -sv2v_cast_D43F7_signed($signed(P[805-:32])) : -sv2v_cast_D43F7_signed($signed(P[611-:32])));
			always @(*) ResNegNF = sv2v_tmp_DB608;
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				case (OutFmt)
					P[773-:2]: ResNegNF = -sv2v_cast_D43F7_signed($signed(P[805-:32]));
					P[579-:2]: ResNegNF = -sv2v_cast_D43F7_signed($signed(P[611-:32]));
					P[449-:2]: ResNegNF = -sv2v_cast_D43F7_signed($signed(P[481-:32]));
					default: ResNegNF = 1'sb0;
				endcase
			end
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				case (OutFmt)
					2'h3: ResNegNF = -sv2v_cast_D43F7_signed($signed(P[1357-:32]));
					2'h1: ResNegNF = -sv2v_cast_D43F7_signed($signed(P[1227-:32]));
					2'h0: ResNegNF = -sv2v_cast_D43F7_signed($signed(P[1097-:32]));
					2'h2: ResNegNF = -sv2v_cast_D43F7_signed($signed(P[967-:32]));
				endcase
			end
		end
	endgenerate
	assign CvtResUf = (($signed(CvtCe) < $signed({{$signed(P[837-:32]) - $clog2($signed(P[805-:32])) {1'b1}}, ResNegNF})) & ~XZero) & ~IntToFp;
	initial _sv2v_0 = 0;
endmodule
module divshiftcalc (
	DivUe,
	DivShiftAmt,
	DivResSubnorm,
	DivSubnormShiftPos
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[837-:32]) + 1:0] DivUe;
	output wire [$signed(P[287-:32]) - 1:0] DivShiftAmt;
	output wire DivResSubnorm;
	output wire DivSubnormShiftPos;
	wire [$signed(P[287-:32]) - 1:0] NormShift;
	wire [$signed(P[287-:32]) - 1:0] DivSubnormShiftAmt;
	wire [$signed(P[837-:32]) + 1:0] DivSubnormShift;
	assign DivResSubnorm = DivUe[$signed(P[837-:32]) + 1] | ~|DivUe[$signed(P[837-:32]) + 1:0];
	function automatic signed [(($signed(P[837-:32]) + 1) >= 0 ? $signed(P[837-:32]) + 2 : 1 - ($signed(P[837-:32]) + 1)) - 1:0] sv2v_cast_A1EFF_signed;
		input reg signed [(($signed(P[837-:32]) + 1) >= 0 ? $signed(P[837-:32]) + 2 : 1 - ($signed(P[837-:32]) + 1)) - 1:0] inp;
		sv2v_cast_A1EFF_signed = inp;
	endfunction
	assign DivSubnormShift = sv2v_cast_A1EFF_signed($signed(P[805-:32])) + DivUe;
	assign DivSubnormShiftPos = ~DivSubnormShift[$signed(P[837-:32]) + 1];
	function automatic signed [$signed(P[287-:32]) - 1:0] sv2v_cast_55618_signed;
		input reg signed [$signed(P[287-:32]) - 1:0] inp;
		sv2v_cast_55618_signed = inp;
	endfunction
	assign NormShift = sv2v_cast_55618_signed($signed(P[805-:32]));
	assign DivSubnormShiftAmt = (DivSubnormShiftPos ? DivSubnormShift[$signed(P[287-:32]) - 1:0] : {$signed(P[287-:32]) {1'sb0}});
	assign DivShiftAmt = (DivResSubnorm ? DivSubnormShiftAmt : NormShift);
endmodule
module flags (
	Xs,
	OutFmt,
	InfIn,
	XInf,
	YInf,
	ZInf,
	NaNIn,
	XSNaN,
	YSNaN,
	ZSNaN,
	XZero,
	YZero,
	FullRe,
	Me,
	Plus1,
	Round,
	Guard,
	Sticky,
	UfPlus1,
	CvtOp,
	ToInt,
	IntToFp,
	Int64,
	Signed,
	CvtCe,
	CvtNegResMsbs,
	DivOp,
	Sqrt,
	FmaOp,
	FmaAs,
	FmaPs,
	DivByZero,
	Overflow,
	Invalid,
	IntInvalid,
	PostProcFlg
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire Xs;
	input wire [$signed(P[707-:32]) - 1:0] OutFmt;
	input wire InfIn;
	input wire XInf;
	input wire YInf;
	input wire ZInf;
	input wire NaNIn;
	input wire XSNaN;
	input wire YSNaN;
	input wire ZSNaN;
	input wire XZero;
	input wire YZero;
	input wire [$signed(P[837-:32]) + 1:0] FullRe;
	input wire [$signed(P[837-:32]) + 1:0] Me;
	input wire Plus1;
	input wire Round;
	input wire Guard;
	input wire Sticky;
	input wire UfPlus1;
	input wire CvtOp;
	input wire ToInt;
	input wire IntToFp;
	input wire Int64;
	input wire Signed;
	input wire [$signed(P[837-:32]):0] CvtCe;
	input wire [1:0] CvtNegResMsbs;
	input wire DivOp;
	input wire Sqrt;
	input wire FmaOp;
	input wire FmaAs;
	input wire FmaPs;
	output wire DivByZero;
	output wire Overflow;
	output wire Invalid;
	output wire IntInvalid;
	output wire [4:0] PostProcFlg;
	wire SigNaN;
	wire Inexact;
	wire FpInexact;
	wire IntInexact;
	wire FmaInvalid;
	wire DivInvalid;
	wire Underflow;
	reg ResExpGteMax;
	wire ShiftGtIntSz;
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk1
			wire [1:1] sv2v_tmp_1480E;
			assign sv2v_tmp_1480E = &FullRe[$signed(P[837-:32]) - 1:0] | FullRe[$signed(P[837-:32])];
			always @(*) ResExpGteMax = sv2v_tmp_1480E;
			assign ShiftGtIntSz = (|FullRe[$signed(P[837-:32]):7] | (FullRe[6] & ~Int64)) | ((|FullRe[4:0] | (FullRe[5] & Int64)) & ((FullRe[5] & ~Int64) | (FullRe[6] & Int64)));
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk1
			wire [1:1] sv2v_tmp_78DAF;
			assign sv2v_tmp_78DAF = (OutFmt ? &FullRe[$signed(P[837-:32]) - 1:0] | FullRe[$signed(P[837-:32])] : &FullRe[$signed(P[643-:32]) - 1:0] | (|FullRe[$signed(P[837-:32]):$signed(P[643-:32])]));
			always @(*) ResExpGteMax = sv2v_tmp_78DAF;
			assign ShiftGtIntSz = (|FullRe[$signed(P[837-:32]):7] | (FullRe[6] & ~Int64)) | ((|FullRe[4:0] | (FullRe[5] & Int64)) & ((FullRe[5] & ~Int64) | (FullRe[6] & Int64)));
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				case (OutFmt)
					P[773-:2]: ResExpGteMax = &FullRe[$signed(P[837-:32]) - 1:0] | FullRe[$signed(P[837-:32])];
					P[579-:2]: ResExpGteMax = &FullRe[$signed(P[643-:32]) - 1:0] | (|FullRe[$signed(P[837-:32]):$signed(P[643-:32])]);
					P[449-:2]: ResExpGteMax = &FullRe[$signed(P[513-:32]) - 1:0] | (|FullRe[$signed(P[837-:32]):$signed(P[513-:32])]);
					default: ResExpGteMax = 1'bx;
				endcase
			end
			assign ShiftGtIntSz = (|FullRe[$signed(P[837-:32]):7] | (FullRe[6] & ~Int64)) | ((|FullRe[4:0] | (FullRe[5] & Int64)) & ((FullRe[5] & ~Int64) | (FullRe[6] & Int64)));
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				case (OutFmt)
					P[1293-:2]: ResExpGteMax = &FullRe[$signed(P[1389-:32]) - 1:0] | FullRe[$signed(P[1389-:32])];
					P[1163-:2]: ResExpGteMax = &FullRe[$signed(P[1259-:32]) - 1:0] | (|FullRe[$signed(P[1389-:32]):$signed(P[1259-:32])]);
					P[1033-:2]: ResExpGteMax = &FullRe[$signed(P[1129-:32]) - 1:0] | (|FullRe[$signed(P[1389-:32]):$signed(P[1129-:32])]);
					P[903-:2]: ResExpGteMax = &FullRe[$signed(P[999-:32]) - 1:0] | (|FullRe[$signed(P[1389-:32]):$signed(P[999-:32])]);
				endcase
			end
			assign ShiftGtIntSz = (|FullRe[$signed(P[1389-:32]):7] | (FullRe[6] & ~Int64)) | ((|FullRe[4:0] | (FullRe[5] & Int64)) & ((FullRe[5] & ~Int64) | (FullRe[6] & Int64)));
		end
	endgenerate
	assign Overflow = (ResExpGteMax & ~FullRe[$signed(P[837-:32]) + 1]) & ~((InfIn | NaNIn) | DivByZero);
	assign Underflow = (((FullRe[$signed(P[837-:32]) + 1] | (FullRe == 0)) | (((FullRe == 1) & (Me == 0)) & ~(UfPlus1 & Guard))) & ((Round | Sticky) | Guard)) & ~(((InfIn | NaNIn) | DivByZero) | Invalid);
	assign FpInexact = (((Sticky | Guard) | Overflow) | Round) & ~(((InfIn | NaNIn) | DivByZero) | Invalid);
	assign IntInexact = ((((CvtCe[$signed(P[837-:32])] & ~XZero) | Sticky) | Round) | Guard) & ~IntInvalid;
	assign Inexact = (ToInt ? IntInexact : FpInexact);
	assign IntInvalid = (((NaNIn | InfIn) | (ShiftGtIntSz & ~FullRe[$signed(P[837-:32]) + 1])) | ((Xs & ~Signed) & ~((CvtCe[$signed(P[837-:32])] | ~|CvtCe) & ~Plus1))) | (CvtNegResMsbs[1] ^ CvtNegResMsbs[0]);
	assign SigNaN = ((XSNaN & ~(IntToFp & CvtOp)) | (YSNaN & ~CvtOp)) | (ZSNaN & FmaOp);
	assign FmaInvalid = (((((XInf | YInf) & ZInf) & (FmaPs ^ FmaAs)) & ~NaNIn) | (XZero & YInf)) | (YZero & XInf);
	assign DivInvalid = (((XInf & YInf) | (XZero & YZero)) & ~Sqrt) | (((Xs & Sqrt) & ~NaNIn) & ~XZero);
	assign Invalid = (SigNaN | (FmaInvalid & FmaOp)) | (DivInvalid & DivOp);
	assign DivByZero = ((YZero & DivOp) & ~Sqrt) & ~((XZero | NaNIn) | InfIn);
	assign PostProcFlg = {Invalid | ((IntInvalid & CvtOp) & ToInt), DivByZero, Overflow & ~(ToInt & CvtOp), Underflow & ~(ToInt & CvtOp), Inexact};
	initial _sv2v_0 = 0;
endmodule
module fmashiftcalc (
	Fmt,
	FmaSe,
	FmaSm,
	FmaSCnt,
	NormSumExp,
	FmaSZero,
	FmaPreResultSubnorm,
	FmaShiftAmt
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[707-:32]) - 1:0] Fmt;
	input wire [$signed(P[837-:32]) + 1:0] FmaSe;
	input wire [$signed(P[255-:32]) - 1:0] FmaSm;
	input wire [$clog2($signed(P[255-:32]) + 1) - 1:0] FmaSCnt;
	output wire [$signed(P[837-:32]) + 1:0] NormSumExp;
	output wire FmaSZero;
	output reg FmaPreResultSubnorm;
	output wire [$clog2($signed(P[255-:32]) + 1) - 1:0] FmaShiftAmt;
	wire [$signed(P[837-:32]) + 1:0] PreNormSumExp;
	reg [$signed(P[837-:32]) + 1:0] BiasCorr;
	assign FmaSZero = ~(|FmaSm);
	function automatic signed [(($signed(P[837-:32]) + 1) >= 0 ? $signed(P[837-:32]) + 2 : 1 - ($signed(P[837-:32]) + 1)) - 1:0] sv2v_cast_A1EFF_signed;
		input reg signed [(($signed(P[837-:32]) + 1) >= 0 ? $signed(P[837-:32]) + 2 : 1 - ($signed(P[837-:32]) + 1)) - 1:0] inp;
		sv2v_cast_A1EFF_signed = inp;
	endfunction
	assign PreNormSumExp = (FmaSe + {{($signed(P[837-:32]) + 2) - $unsigned($clog2($signed(P[255-:32]) + 1)) {1'b1}}, ~FmaSCnt}) + sv2v_cast_A1EFF_signed($signed(P[805-:32]) + 4);
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk1
			assign NormSumExp = PreNormSumExp;
			wire [(($signed(P[837-:32]) + 1) >= 0 ? $signed(P[837-:32]) + 2 : 1 - ($signed(P[837-:32]) + 1)):1] sv2v_tmp_591EA;
			assign sv2v_tmp_591EA = 1'sb0;
			always @(*) BiasCorr = sv2v_tmp_591EA;
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk1
			wire [(($signed(P[837-:32]) + 1) >= 0 ? $signed(P[837-:32]) + 2 : 1 - ($signed(P[837-:32]) + 1)):1] sv2v_tmp_1001D;
			assign sv2v_tmp_1001D = (Fmt ? sv2v_cast_A1EFF_signed(0) : sv2v_cast_A1EFF_signed($signed(P[577-:32]) - $signed(P[771-:32])));
			always @(*) BiasCorr = sv2v_tmp_1001D;
			assign NormSumExp = PreNormSumExp + BiasCorr;
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					P[773-:2]: BiasCorr = 1'sb0;
					P[579-:2]: BiasCorr = sv2v_cast_A1EFF_signed($signed(P[577-:32]) - $signed(P[771-:32]));
					P[449-:2]: BiasCorr = sv2v_cast_A1EFF_signed($signed(P[447-:32]) - $signed(P[771-:32]));
					default: BiasCorr = 1'sbx;
				endcase
			end
			assign NormSumExp = PreNormSumExp + BiasCorr;
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					2'h3: BiasCorr = 1'sb0;
					2'h1: BiasCorr = sv2v_cast_A1EFF_signed($signed(P[1195-:32]) - $signed(P[1325-:32]));
					2'h0: BiasCorr = sv2v_cast_A1EFF_signed($signed(P[1065-:32]) - $signed(P[1325-:32]));
					2'h2: BiasCorr = sv2v_cast_A1EFF_signed($signed(P[935-:32]) - $signed(P[1325-:32]));
				endcase
			end
			assign NormSumExp = PreNormSumExp + BiasCorr;
		end
		if ($signed(P[739-:32]) == 1) begin : genblk2
			wire Sum0LEZ;
			wire Sum0GEFL;
			assign Sum0LEZ = PreNormSumExp[$signed(P[837-:32]) + 1] | ~|PreNormSumExp;
			assign Sum0GEFL = $signed(PreNormSumExp) >= $signed(sv2v_cast_A1EFF_signed(-($signed(P[805-:32]) + 1)));
			wire [1:1] sv2v_tmp_7BA83;
			assign sv2v_tmp_7BA83 = Sum0LEZ & Sum0GEFL;
			always @(*) FmaPreResultSubnorm = sv2v_tmp_7BA83;
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk2
			wire Sum0LEZ;
			wire Sum0GEFL;
			wire Sum1LEZ;
			wire Sum1GEFL;
			assign Sum0LEZ = PreNormSumExp[$signed(P[837-:32]) + 1] | ~|PreNormSumExp;
			assign Sum0GEFL = $signed(PreNormSumExp) >= $signed(sv2v_cast_A1EFF_signed(-($signed(P[805-:32]) + 1)));
			assign Sum1LEZ = $signed(PreNormSumExp) <= $signed(sv2v_cast_A1EFF_signed($signed(P[771-:32]) - $signed(P[577-:32])));
			assign Sum1GEFL = ($signed(PreNormSumExp) >= $signed(sv2v_cast_A1EFF_signed(($signed(P[771-:32]) - ($signed(P[611-:32]) + 1)) - $signed(P[577-:32])))) | ~|PreNormSumExp;
			wire [1:1] sv2v_tmp_6615D;
			assign sv2v_tmp_6615D = (Fmt ? Sum0LEZ : Sum1LEZ) & (Fmt ? Sum0GEFL : Sum1GEFL);
			always @(*) FmaPreResultSubnorm = sv2v_tmp_6615D;
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk2
			wire Sum0LEZ;
			wire Sum0GEFL;
			wire Sum1LEZ;
			wire Sum1GEFL;
			wire Sum2LEZ;
			wire Sum2GEFL;
			assign Sum0LEZ = PreNormSumExp[$signed(P[837-:32]) + 1] | ~|PreNormSumExp;
			assign Sum0GEFL = $signed(PreNormSumExp) >= $signed(sv2v_cast_A1EFF_signed(-($signed(P[805-:32]) + 1)));
			assign Sum1LEZ = $signed(PreNormSumExp) <= $signed(sv2v_cast_A1EFF_signed($signed(P[771-:32]) - $signed(P[577-:32])));
			assign Sum1GEFL = ($signed(PreNormSumExp) >= $signed(sv2v_cast_A1EFF_signed(($signed(P[771-:32]) - ($signed(P[611-:32]) + 1)) - $signed(P[577-:32])))) | ~|PreNormSumExp;
			assign Sum2LEZ = $signed(PreNormSumExp) <= $signed(sv2v_cast_A1EFF_signed($signed(P[771-:32]) - $signed(P[447-:32])));
			assign Sum2GEFL = ($signed(PreNormSumExp) >= $signed(sv2v_cast_A1EFF_signed(($signed(P[771-:32]) - ($signed(P[481-:32]) + 1)) - $signed(P[447-:32])))) | ~|PreNormSumExp;
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					P[773-:2]: FmaPreResultSubnorm = Sum0LEZ & Sum0GEFL;
					P[579-:2]: FmaPreResultSubnorm = Sum1LEZ & Sum1GEFL;
					P[449-:2]: FmaPreResultSubnorm = Sum2LEZ & Sum2GEFL;
					default: FmaPreResultSubnorm = 1'bx;
				endcase
			end
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk2
			wire Sum0LEZ;
			wire Sum0GEFL;
			wire Sum1LEZ;
			wire Sum1GEFL;
			wire Sum2LEZ;
			wire Sum2GEFL;
			wire Sum3LEZ;
			wire Sum3GEFL;
			assign Sum0LEZ = PreNormSumExp[$signed(P[837-:32]) + 1] | ~|PreNormSumExp;
			assign Sum0GEFL = $signed(PreNormSumExp) >= $signed(sv2v_cast_A1EFF_signed(-($signed(P[805-:32]) + 1)));
			assign Sum1LEZ = $signed(PreNormSumExp) <= $signed(sv2v_cast_A1EFF_signed($signed(P[771-:32]) - $signed(P[1195-:32])));
			assign Sum1GEFL = ($signed(PreNormSumExp) >= $signed(sv2v_cast_A1EFF_signed(($signed(P[771-:32]) - ($signed(P[1227-:32]) + 1)) - $signed(P[1195-:32])))) | ~|PreNormSumExp;
			assign Sum2LEZ = $signed(PreNormSumExp) <= $signed(sv2v_cast_A1EFF_signed($signed(P[771-:32]) - $signed(P[1065-:32])));
			assign Sum2GEFL = ($signed(PreNormSumExp) >= $signed(sv2v_cast_A1EFF_signed(($signed(P[771-:32]) - ($signed(P[1097-:32]) + 1)) - $signed(P[1065-:32])))) | ~|PreNormSumExp;
			assign Sum3LEZ = $signed(PreNormSumExp) <= $signed(sv2v_cast_A1EFF_signed($signed(P[771-:32]) - $signed(P[935-:32])));
			assign Sum3GEFL = ($signed(PreNormSumExp) >= $signed(sv2v_cast_A1EFF_signed(($signed(P[771-:32]) - ($signed(P[967-:32]) + 1)) - $signed(P[935-:32])))) | ~|PreNormSumExp;
			always @(*) begin
				if (_sv2v_0)
					;
				case (Fmt)
					2'h3: FmaPreResultSubnorm = Sum0LEZ & Sum0GEFL;
					2'h1: FmaPreResultSubnorm = Sum1LEZ & Sum1GEFL;
					2'h0: FmaPreResultSubnorm = Sum2LEZ & Sum2GEFL;
					2'h2: FmaPreResultSubnorm = Sum3LEZ & Sum3GEFL;
				endcase
			end
		end
	endgenerate
	function automatic signed [$clog2($signed(P[255-:32]) - 1) - 1:0] sv2v_cast_E062E_signed;
		input reg signed [$clog2($signed(P[255-:32]) - 1) - 1:0] inp;
		sv2v_cast_E062E_signed = inp;
	endfunction
	assign FmaShiftAmt = (FmaPreResultSubnorm ? (FmaSe[$clog2($signed(P[255-:32]) - 1) - 1:0] + sv2v_cast_E062E_signed($signed(P[805-:32]) + 3)) + BiasCorr[$clog2($signed(P[255-:32]) - 1) - 1:0] : FmaSCnt + 1);
	initial _sv2v_0 = 0;
endmodule
module negateintres (
	Signed,
	Int64,
	Plus1,
	Xs,
	Shifted,
	CvtNegResMsbs,
	CvtNegRes
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire Signed;
	input wire Int64;
	input wire Plus1;
	input wire Xs;
	input wire [$signed(P[319-:32]) - 1:0] Shifted;
	output wire [1:0] CvtNegResMsbs;
	output wire [$signed(P[4216-:32]) + 1:0] CvtNegRes;
	wire [$signed(P[4216-:32]) + 1:0] CvtPreRes;
	wire [2:0] CvtNegResMsbs3;
	assign CvtPreRes = {2'b00, Shifted[$signed(P[319-:32]) - 1:$signed(P[319-:32]) - $signed(P[4216-:32])]} + {{$signed(P[4216-:32]) + 1 {1'b0}}, Plus1};
	mux2 #(.WIDTH($signed(P[4216-:32]) + 2)) resmux(
		.d0(CvtPreRes),
		.d1(-CvtPreRes),
		.s(Xs),
		.y(CvtNegRes)
	);
	mux2 #(.WIDTH(3)) msb3mux(
		.d0(CvtNegRes[33:31]),
		.d1(CvtNegRes[$signed(P[4216-:32]) + 1:$signed(P[4216-:32]) - 1]),
		.s(Int64),
		.y(CvtNegResMsbs3)
	);
	mux2 #(.WIDTH(2)) msb2mux(
		.d0(CvtNegResMsbs3[2:1]),
		.d1(CvtNegResMsbs3[1:0]),
		.s(Signed),
		.y(CvtNegResMsbs)
	);
endmodule
module normshift (
	ShiftAmt,
	ShiftIn,
	Shifted
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[287-:32]) - 1:0] ShiftAmt;
	input wire [$signed(P[319-:32]) - 1:0] ShiftIn;
	output wire [$signed(P[319-:32]) - 1:0] Shifted;
	assign Shifted = ShiftIn << ShiftAmt;
endmodule
module postprocess (
	Xs,
	Ys,
	Xm,
	Ym,
	Zm,
	Frm,
	Fmt,
	OpCtrl,
	XZero,
	YZero,
	XInf,
	YInf,
	ZInf,
	XNaN,
	YNaN,
	ZNaN,
	XSNaN,
	YSNaN,
	ZSNaN,
	PostProcSel,
	FmaAs,
	FmaPs,
	FmaSs,
	FmaSe,
	FmaSm,
	FmaASticky,
	FmaSCnt,
	DivSticky,
	DivUe,
	DivUm,
	CvtCs,
	CvtCe,
	CvtResSubnormUf,
	CvtShiftAmt,
	ToInt,
	Zfa,
	CvtLzcIn,
	IntZero,
	PostProcRes,
	PostProcFlg,
	FCvtIntRes
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire Xs;
	input wire Ys;
	input wire [$signed(P[805-:32]):0] Xm;
	input wire [$signed(P[805-:32]):0] Ym;
	input wire [$signed(P[805-:32]):0] Zm;
	input wire [2:0] Frm;
	input wire [$signed(P[707-:32]) - 1:0] Fmt;
	input wire [2:0] OpCtrl;
	input wire XZero;
	input wire YZero;
	input wire XInf;
	input wire YInf;
	input wire ZInf;
	input wire XNaN;
	input wire YNaN;
	input wire ZNaN;
	input wire XSNaN;
	input wire YSNaN;
	input wire ZSNaN;
	input wire [1:0] PostProcSel;
	input wire FmaAs;
	input wire FmaPs;
	input wire FmaSs;
	input wire [$signed(P[837-:32]) + 1:0] FmaSe;
	input wire [$signed(P[255-:32]) - 1:0] FmaSm;
	input wire FmaASticky;
	input wire [$clog2($signed(P[255-:32]) + 1) - 1:0] FmaSCnt;
	input wire DivSticky;
	input wire [$signed(P[837-:32]) + 1:0] DivUe;
	input wire [$signed(P[95-:32]):0] DivUm;
	input wire CvtCs;
	input wire [$signed(P[837-:32]):0] CvtCe;
	input wire CvtResSubnormUf;
	input wire [$signed(P[351-:32]) - 1:0] CvtShiftAmt;
	input wire ToInt;
	input wire Zfa;
	input wire [$signed(P[415-:32]) - 1:0] CvtLzcIn;
	input wire IntZero;
	output wire [$signed(P[901-:32]) - 1:0] PostProcRes;
	output wire [4:0] PostProcFlg;
	output wire [$signed(P[4216-:32]) - 1:0] FCvtIntRes;
	wire Rs;
	wire [$signed(P[805-:32]) - 1:0] Rf;
	wire [$signed(P[837-:32]) - 1:0] Re;
	wire Ms;
	wire [$signed(P[319-:32]) - 1:0] Mf;
	wire [$signed(P[837-:32]) + 1:0] Me;
	wire [$signed(P[837-:32]) + 1:0] FullRe;
	wire UfPlus1;
	reg [$signed(P[287-:32]) - 1:0] ShiftAmt;
	reg [$signed(P[319-:32]) - 1:0] ShiftIn;
	wire [$signed(P[319-:32]) - 1:0] Shifted;
	wire Plus1;
	wire Overflow;
	wire Invalid;
	wire Guard;
	wire Round;
	wire Sticky;
	wire [$signed(P[707-:32]) - 1:0] OutFmt;
	wire [$signed(P[837-:32]) + 1:0] FmaMe;
	wire FmaSZero;
	wire [$signed(P[837-:32]) + 1:0] NormSumExp;
	wire FmaPreResultSubnorm;
	wire [$clog2($signed(P[255-:32]) + 1) - 1:0] FmaShiftAmt;
	wire [$signed(P[287-:32]) - 1:0] DivShiftAmt;
	wire [$signed(P[837-:32]) + 1:0] Ue;
	wire DivByZero;
	wire DivResSubnorm;
	wire DivSubnormShiftPos;
	wire [$signed(P[415-:32]) + $signed(P[805-:32]):0] CvtShiftIn;
	wire [1:0] CvtNegResMsbs;
	wire [$signed(P[4216-:32]) + 1:0] CvtNegRes;
	wire CvtResUf;
	wire IntInvalid;
	wire Mult;
	wire Sqrt;
	wire Int64;
	wire Signed;
	wire IntToFp;
	wire CvtOp;
	wire FmaOp;
	wire DivOp;
	wire InfIn;
	wire NaNIn;
	assign Signed = OpCtrl[0];
	assign Int64 = OpCtrl[1];
	assign IntToFp = OpCtrl[2];
	assign Mult = (OpCtrl[2] & ~OpCtrl[1]) & ~OpCtrl[0];
	assign CvtOp = PostProcSel == 2'b00;
	assign FmaOp = PostProcSel == 2'b10;
	assign DivOp = PostProcSel == 2'b01;
	assign Sqrt = OpCtrl[0];
	assign InfIn = (XInf | YInf) | ZInf;
	assign NaNIn = (XNaN | YNaN) | ZNaN;
	generate
		if ($signed(P[739-:32]) == 2) begin : genblk1
			assign OutFmt = (IntToFp | ~CvtOp ? Fmt : OpCtrl[1:0] == P[773-:2]);
		end
		else if (($signed(P[739-:32]) == 3) | ($signed(P[739-:32]) == 4)) begin : genblk1
			assign OutFmt = (IntToFp | ~CvtOp ? Fmt : OpCtrl[1:0]);
		end
		else begin : genblk1
			assign OutFmt = 0;
		end
	endgenerate
	cvtshiftcalc #(.P(P)) cvtshiftcalc(
		.ToInt(ToInt),
		.CvtCe(CvtCe),
		.CvtResSubnormUf(CvtResSubnormUf),
		.Xm(Xm),
		.CvtLzcIn(CvtLzcIn),
		.XZero(XZero),
		.IntToFp(IntToFp),
		.OutFmt(OutFmt),
		.CvtResUf(CvtResUf),
		.CvtShiftIn(CvtShiftIn)
	);
	fmashiftcalc #(.P(P)) fmashiftcalc(
		.FmaSCnt(FmaSCnt),
		.Fmt(Fmt),
		.NormSumExp(NormSumExp),
		.FmaSe(FmaSe),
		.FmaSm(FmaSm),
		.FmaSZero(FmaSZero),
		.FmaPreResultSubnorm(FmaPreResultSubnorm),
		.FmaShiftAmt(FmaShiftAmt)
	);
	divshiftcalc #(.P(P)) divshiftcalc(
		.DivUe(DivUe),
		.DivResSubnorm(DivResSubnorm),
		.DivSubnormShiftPos(DivSubnormShiftPos),
		.DivShiftAmt(DivShiftAmt)
	);
	always @(*) begin
		if (_sv2v_0)
			;
		case (PostProcSel)
			2'b10: begin
				ShiftAmt = {{$signed(P[287-:32]) - $clog2($signed(P[255-:32]) - 1) {1'b0}}, FmaShiftAmt};
				ShiftIn = {2'b00, FmaSm, {$signed(P[319-:32]) - ($signed(P[255-:32]) + 2) {1'b0}}};
			end
			2'b00: begin
				ShiftAmt = {{$signed(P[287-:32]) - $clog2($signed(P[415-:32]) + 1) {1'b0}}, CvtShiftAmt};
				ShiftIn = {CvtShiftIn, {$signed(P[319-:32]) - (($signed(P[415-:32]) + $signed(P[805-:32])) + 1) {1'b0}}};
			end
			2'b01: begin
				ShiftAmt = DivShiftAmt;
				ShiftIn = {{$signed(P[805-:32]) {1'b0}}, DivUm, {$signed(P[319-:32]) - (($signed(P[95-:32]) + 1) + $signed(P[805-:32])) {1'b0}}};
			end
			default: begin
				ShiftAmt = {$signed(P[287-:32]) {1'bx}};
				ShiftIn = {$signed(P[319-:32]) {1'bx}};
			end
		endcase
	end
	normshift #(.P(P)) normshift(
		.ShiftIn(ShiftIn),
		.ShiftAmt(ShiftAmt),
		.Shifted(Shifted)
	);
	shiftcorrection #(.P(P)) shiftcorrection(
		.FmaOp(FmaOp),
		.FmaPreResultSubnorm(FmaPreResultSubnorm),
		.NormSumExp(NormSumExp),
		.DivResSubnorm(DivResSubnorm),
		.DivSubnormShiftPos(DivSubnormShiftPos),
		.DivOp(DivOp),
		.DivUe(DivUe),
		.Ue(Ue),
		.FmaSZero(FmaSZero),
		.Shifted(Shifted),
		.FmaMe(FmaMe),
		.Mf(Mf)
	);
	roundsign roundsign(
		.FmaOp(FmaOp),
		.DivOp(DivOp),
		.CvtOp(CvtOp),
		.Sqrt(Sqrt),
		.FmaSs(FmaSs),
		.Xs(Xs),
		.Ys(Ys),
		.CvtCs(CvtCs),
		.Ms(Ms)
	);
	round #(.P(P)) round(
		.OutFmt(OutFmt),
		.Frm(Frm),
		.FmaASticky(FmaASticky),
		.Plus1(Plus1),
		.PostProcSel(PostProcSel),
		.CvtCe(CvtCe),
		.Ue(Ue),
		.Ms(Ms),
		.FmaMe(FmaMe),
		.FmaOp(FmaOp),
		.CvtOp(CvtOp),
		.CvtResSubnormUf(CvtResSubnormUf),
		.Mf(Mf),
		.ToInt(ToInt),
		.CvtResUf(CvtResUf),
		.DivSticky(DivSticky),
		.DivOp(DivOp),
		.UfPlus1(UfPlus1),
		.FullRe(FullRe),
		.Rf(Rf),
		.Re(Re),
		.Sticky(Sticky),
		.Round(Round),
		.Guard(Guard),
		.Me(Me)
	);
	resultsign resultsign(
		.Frm(Frm),
		.FmaPs(FmaPs),
		.FmaAs(FmaAs),
		.Round(Round),
		.Sticky(Sticky),
		.Guard(Guard),
		.FmaOp(FmaOp),
		.ZInf(ZInf),
		.InfIn(InfIn),
		.FmaSZero(FmaSZero),
		.Mult(Mult),
		.Ms(Ms),
		.Rs(Rs)
	);
	flags #(.P(P)) flags(
		.XSNaN(XSNaN),
		.YSNaN(YSNaN),
		.ZSNaN(ZSNaN),
		.XInf(XInf),
		.YInf(YInf),
		.ZInf(ZInf),
		.InfIn(InfIn),
		.XZero(XZero),
		.YZero(YZero),
		.Xs(Xs),
		.Sqrt(Sqrt),
		.ToInt(ToInt),
		.IntToFp(IntToFp),
		.Int64(Int64),
		.Signed(Signed),
		.OutFmt(OutFmt),
		.CvtCe(CvtCe),
		.NaNIn(NaNIn),
		.FmaAs(FmaAs),
		.FmaPs(FmaPs),
		.Round(Round),
		.IntInvalid(IntInvalid),
		.DivByZero(DivByZero),
		.Guard(Guard),
		.Sticky(Sticky),
		.UfPlus1(UfPlus1),
		.CvtOp(CvtOp),
		.DivOp(DivOp),
		.FmaOp(FmaOp),
		.FullRe(FullRe),
		.Plus1(Plus1),
		.Me(Me),
		.CvtNegResMsbs(CvtNegResMsbs),
		.Invalid(Invalid),
		.Overflow(Overflow),
		.PostProcFlg(PostProcFlg)
	);
	negateintres #(.P(P)) negateintres(
		.Xs(Xs),
		.Shifted(Shifted),
		.Signed(Signed),
		.Int64(Int64),
		.Plus1(Plus1),
		.CvtNegResMsbs(CvtNegResMsbs),
		.CvtNegRes(CvtNegRes)
	);
	specialcase #(.P(P)) specialcase(
		.Xs(Xs),
		.Xm(Xm),
		.Ym(Ym),
		.Zm(Zm),
		.XZero(XZero),
		.IntInvalid(IntInvalid),
		.IntZero(IntZero),
		.Frm(Frm),
		.OutFmt(OutFmt),
		.XNaN(XNaN),
		.YNaN(YNaN),
		.ZNaN(ZNaN),
		.CvtResUf(CvtResUf),
		.NaNIn(NaNIn),
		.IntToFp(IntToFp),
		.Int64(Int64),
		.Signed(Signed),
		.Zfa(Zfa),
		.CvtOp(CvtOp),
		.FmaOp(FmaOp),
		.Plus1(Plus1),
		.Invalid(Invalid),
		.Overflow(Overflow),
		.InfIn(InfIn),
		.CvtNegRes(CvtNegRes),
		.XInf(XInf),
		.YInf(YInf),
		.DivOp(DivOp),
		.DivByZero(DivByZero),
		.FullRe(FullRe),
		.CvtCe(CvtCe),
		.Rs(Rs),
		.Re(Re),
		.Rf(Rf),
		.PostProcRes(PostProcRes),
		.FCvtIntRes(FCvtIntRes)
	);
	initial _sv2v_0 = 0;
endmodule
module resultsign (
	Frm,
	FmaOp,
	Mult,
	ZInf,
	InfIn,
	FmaSZero,
	Ms,
	FmaPs,
	FmaAs,
	Guard,
	Round,
	Sticky,
	Rs
);
	reg _sv2v_0;
	input wire [2:0] Frm;
	input wire FmaOp;
	input wire Mult;
	input wire ZInf;
	input wire InfIn;
	input wire FmaSZero;
	input wire Ms;
	input wire FmaPs;
	input wire FmaAs;
	input wire Guard;
	input wire Round;
	input wire Sticky;
	output reg Rs;
	wire Zeros;
	wire Infs;
	assign Zeros = (((FmaPs ^ FmaAs) & ~((Round | Guard) | Sticky)) & ~Mult ? Frm[1:0] == 2'b10 : FmaPs);
	assign Infs = (ZInf ? FmaAs : FmaPs);
	always @(*) begin
		if (_sv2v_0)
			;
		if (InfIn & FmaOp)
			Rs = Infs;
		else if (FmaSZero & FmaOp)
			Rs = Zeros;
		else
			Rs = Ms;
	end
	initial _sv2v_0 = 0;
endmodule
module round (
	OutFmt,
	Frm,
	PostProcSel,
	Ms,
	Mf,
	FmaOp,
	FmaMe,
	FmaASticky,
	DivOp,
	DivSticky,
	Ue,
	CvtOp,
	ToInt,
	CvtResSubnormUf,
	CvtResUf,
	CvtCe,
	Me,
	UfPlus1,
	FullRe,
	Re,
	Rf,
	Sticky,
	Plus1,
	Round,
	Guard
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[707-:32]) - 1:0] OutFmt;
	input wire [2:0] Frm;
	input wire [1:0] PostProcSel;
	input wire Ms;
	input wire [$signed(P[319-:32]) - 1:0] Mf;
	input wire FmaOp;
	input wire [$signed(P[837-:32]) + 1:0] FmaMe;
	input wire FmaASticky;
	input wire DivOp;
	input wire DivSticky;
	input wire [$signed(P[837-:32]) + 1:0] Ue;
	input wire CvtOp;
	input wire ToInt;
	input wire CvtResSubnormUf;
	input wire CvtResUf;
	input wire [$signed(P[837-:32]):0] CvtCe;
	output reg [$signed(P[837-:32]) + 1:0] Me;
	output wire UfPlus1;
	output wire [$signed(P[837-:32]) + 1:0] FullRe;
	output wire [$signed(P[837-:32]) - 1:0] Re;
	output wire [$signed(P[805-:32]) - 1:0] Rf;
	output wire Sticky;
	output wire Plus1;
	output wire Round;
	output wire Guard;
	reg UfCalcPlus1;
	wire NormSticky;
	wire [$signed(P[805-:32]) - 1:0] RoundFrac;
	wire FpRes;
	wire IntRes;
	reg FpGuard;
	reg FpRound;
	reg FpLsbRes;
	wire LsbRes;
	reg CalcPlus1;
	wire FpPlus1;
	wire [$signed(P[901-:32]):0] RoundAdd;
	wire CvtToInt;
	localparam XLENPOS = ($signed(P[4216-:32]) > $signed(P[805-:32]) ? 1 : ($signed(P[4216-:32]) > $signed(P[611-:32]) ? 2 : 3));
	assign IntRes = ToInt;
	assign FpRes = ~IntRes;
	assign CvtToInt = ToInt;
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk1
			if (XLENPOS == 1) begin : genblk1
				assign NormSticky = (|Mf[($signed(P[319-:32]) - $signed(P[805-:32])) - 2:($signed(P[319-:32]) - $signed(P[4216-:32])) - 1] & FpRes) | (|Mf[($signed(P[319-:32]) - $signed(P[4216-:32])) - 2:0]);
			end
			if (XLENPOS == 2) begin : genblk2
				assign NormSticky = (|Mf[($signed(P[319-:32]) - $signed(P[4216-:32])) - 2:($signed(P[319-:32]) - $signed(P[805-:32])) - 1] & IntRes) | (|Mf[($signed(P[319-:32]) - $signed(P[805-:32])) - 2:0]);
			end
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk1
			if (XLENPOS == 1) begin : genblk1
				assign NormSticky = (((|Mf[($signed(P[319-:32]) - $signed(P[611-:32])) - 2:($signed(P[319-:32]) - $signed(P[805-:32])) - 1] & FpRes) & ~OutFmt) | (|Mf[($signed(P[319-:32]) - $signed(P[805-:32])) - 2:($signed(P[319-:32]) - $signed(P[4216-:32])) - 1] & FpRes)) | (|Mf[($signed(P[319-:32]) - $signed(P[4216-:32])) - 2:0]);
			end
			if (XLENPOS == 2) begin : genblk2
				assign NormSticky = (((|Mf[($signed(P[319-:32]) - $signed(P[611-:32])) - 2:($signed(P[319-:32]) - $signed(P[4216-:32])) - 1] & FpRes) & ~OutFmt) | (|Mf[($signed(P[319-:32]) - $signed(P[4216-:32])) - 2:($signed(P[319-:32]) - $signed(P[805-:32])) - 1] & (IntRes | ~OutFmt))) | (|Mf[($signed(P[319-:32]) - $signed(P[805-:32])) - 2:0]);
			end
			if (XLENPOS == 3) begin : genblk3
				assign NormSticky = ((|Mf[($signed(P[319-:32]) - $signed(P[4216-:32])) - 2:($signed(P[319-:32]) - $signed(P[611-:32])) - 1] & IntRes) | (|Mf[($signed(P[319-:32]) - $signed(P[611-:32])) - 2:($signed(P[319-:32]) - $signed(P[805-:32])) - 1] & (~OutFmt | IntRes))) | (|Mf[($signed(P[319-:32]) - $signed(P[805-:32])) - 2:0]);
			end
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk1
			if (XLENPOS == 1) begin : genblk1
				assign NormSticky = ((((|Mf[($signed(P[319-:32]) - $signed(P[481-:32])) - 2:($signed(P[319-:32]) - $signed(P[611-:32])) - 1] & FpRes) & (OutFmt == P[449-:2])) | ((|Mf[($signed(P[319-:32]) - $signed(P[611-:32])) - 2:($signed(P[319-:32]) - $signed(P[805-:32])) - 1] & FpRes) & ~(OutFmt == P[773-:2]))) | (|Mf[($signed(P[319-:32]) - $signed(P[805-:32])) - 2:($signed(P[319-:32]) - $signed(P[4216-:32])) - 1] & FpRes)) | (|Mf[($signed(P[319-:32]) - $signed(P[4216-:32])) - 2:0]);
			end
			if (XLENPOS == 2) begin : genblk2
				assign NormSticky = ((((|Mf[($signed(P[319-:32]) - $signed(P[481-:32])) - 2:($signed(P[319-:32]) - $signed(P[611-:32])) - 1] & FpRes) & (OutFmt == P[449-:2])) | ((|Mf[($signed(P[319-:32]) - $signed(P[611-:32])) - 2:($signed(P[319-:32]) - $signed(P[4216-:32])) - 1] & FpRes) & ~(OutFmt == P[773-:2]))) | (|Mf[($signed(P[319-:32]) - $signed(P[4216-:32])) - 2:($signed(P[319-:32]) - $signed(P[805-:32])) - 1] & (IntRes | ~(OutFmt == P[773-:2])))) | (|Mf[($signed(P[319-:32]) - $signed(P[805-:32])) - 2:0]);
			end
			if (XLENPOS == 3) begin : genblk3
				assign NormSticky = ((((|Mf[($signed(P[319-:32]) - $signed(P[481-:32])) - 2:($signed(P[319-:32]) - $signed(P[4216-:32])) - 1] & FpRes) & (OutFmt == P[449-:2])) | (|Mf[($signed(P[319-:32]) - $signed(P[4216-:32])) - 2:($signed(P[319-:32]) - $signed(P[611-:32])) - 1] & ((OutFmt == P[449-:2]) | IntRes))) | (|Mf[($signed(P[319-:32]) - $signed(P[611-:32])) - 2:($signed(P[319-:32]) - $signed(P[805-:32])) - 1] & (~(OutFmt == P[773-:2]) | IntRes))) | (|Mf[($signed(P[319-:32]) - $signed(P[805-:32])) - 2:0]);
			end
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk1
			if (XLENPOS == 2) begin : genblk1
				assign NormSticky = (((((|Mf[($signed(P[319-:32]) - $signed(P[967-:32])) - 2:($signed(P[319-:32]) - $signed(P[1097-:32])) - 1] & FpRes) & (OutFmt == P[903-:2])) | ((|Mf[($signed(P[319-:32]) - $signed(P[1097-:32])) - 2:($signed(P[319-:32]) - $signed(P[1227-:32])) - 1] & FpRes) & ((OutFmt == P[1033-:2]) | (OutFmt == P[903-:2])))) | ((|Mf[($signed(P[319-:32]) - $signed(P[1227-:32])) - 2:($signed(P[319-:32]) - $signed(P[4216-:32])) - 1] & FpRes) & ~(OutFmt == P[1293-:2]))) | (|Mf[($signed(P[319-:32]) - $signed(P[4216-:32])) - 2:($signed(P[319-:32]) - $signed(P[1357-:32])) - 1] & (~(OutFmt == P[1293-:2]) | IntRes))) | (|Mf[($signed(P[319-:32]) - $signed(P[1357-:32])) - 2:0]);
			end
			if (XLENPOS == 3) begin : genblk2
				assign NormSticky = (((((|Mf[($signed(P[319-:32]) - $signed(P[967-:32])) - 2:($signed(P[319-:32]) - $signed(P[1097-:32])) - 1] & FpRes) & (OutFmt == P[903-:2])) | ((|Mf[($signed(P[319-:32]) - $signed(P[1097-:32])) - 2:($signed(P[319-:32]) - $signed(P[4216-:32])) - 1] & FpRes) & ((OutFmt == P[1033-:2]) | (OutFmt == P[903-:2])))) | (|Mf[($signed(P[319-:32]) - $signed(P[4216-:32])) - 2:($signed(P[319-:32]) - $signed(P[1227-:32])) - 1] & (((OutFmt == P[1033-:2]) | (OutFmt == P[903-:2])) | IntRes))) | (|Mf[($signed(P[319-:32]) - $signed(P[1227-:32])) - 2:($signed(P[319-:32]) - $signed(P[1357-:32])) - 1] & (~(OutFmt == P[1293-:2]) | IntRes))) | (|Mf[($signed(P[319-:32]) - $signed(P[1357-:32])) - 2:0]);
			end
		end
	endgenerate
	assign Sticky = ((((FmaASticky & FmaOp) | NormSticky) | (CvtResUf & CvtOp)) | (FmaMe[$signed(P[837-:32]) + 1] & FmaOp)) | (DivSticky & DivOp);
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk2
			wire [1:1] sv2v_tmp_A50F1;
			assign sv2v_tmp_A50F1 = Mf[($signed(P[319-:32]) - $signed(P[805-:32])) - 1];
			always @(*) FpGuard = sv2v_tmp_A50F1;
			wire [1:1] sv2v_tmp_16C3B;
			assign sv2v_tmp_16C3B = Mf[$signed(P[319-:32]) - $signed(P[805-:32])];
			always @(*) FpLsbRes = sv2v_tmp_16C3B;
			wire [1:1] sv2v_tmp_25B95;
			assign sv2v_tmp_25B95 = Mf[($signed(P[319-:32]) - $signed(P[805-:32])) - 2];
			always @(*) FpRound = sv2v_tmp_25B95;
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk2
			wire [1:1] sv2v_tmp_4941A;
			assign sv2v_tmp_4941A = (OutFmt ? Mf[($signed(P[319-:32]) - $signed(P[805-:32])) - 1] : Mf[($signed(P[319-:32]) - $signed(P[611-:32])) - 1]);
			always @(*) FpGuard = sv2v_tmp_4941A;
			wire [1:1] sv2v_tmp_17D79;
			assign sv2v_tmp_17D79 = (OutFmt ? Mf[$signed(P[319-:32]) - $signed(P[805-:32])] : Mf[$signed(P[319-:32]) - $signed(P[611-:32])]);
			always @(*) FpLsbRes = sv2v_tmp_17D79;
			wire [1:1] sv2v_tmp_4681D;
			assign sv2v_tmp_4681D = (OutFmt ? Mf[($signed(P[319-:32]) - $signed(P[805-:32])) - 2] : Mf[($signed(P[319-:32]) - $signed(P[611-:32])) - 2]);
			always @(*) FpRound = sv2v_tmp_4681D;
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk2
			always @(*) begin
				if (_sv2v_0)
					;
				case (OutFmt)
					P[773-:2]: begin
						FpGuard = Mf[($signed(P[319-:32]) - $signed(P[805-:32])) - 1];
						FpLsbRes = Mf[$signed(P[319-:32]) - $signed(P[805-:32])];
						FpRound = Mf[($signed(P[319-:32]) - $signed(P[805-:32])) - 2];
					end
					P[579-:2]: begin
						FpGuard = Mf[($signed(P[319-:32]) - $signed(P[611-:32])) - 1];
						FpLsbRes = Mf[$signed(P[319-:32]) - $signed(P[611-:32])];
						FpRound = Mf[($signed(P[319-:32]) - $signed(P[611-:32])) - 2];
					end
					P[449-:2]: begin
						FpGuard = Mf[($signed(P[319-:32]) - $signed(P[481-:32])) - 1];
						FpLsbRes = Mf[$signed(P[319-:32]) - $signed(P[481-:32])];
						FpRound = Mf[($signed(P[319-:32]) - $signed(P[481-:32])) - 2];
					end
					default: begin
						FpGuard = 1'bx;
						FpLsbRes = 1'bx;
						FpRound = 1'bx;
					end
				endcase
			end
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk2
			always @(*) begin
				if (_sv2v_0)
					;
				case (OutFmt)
					2'h3: begin
						FpGuard = Mf[($signed(P[319-:32]) - $signed(P[1357-:32])) - 1];
						FpLsbRes = Mf[$signed(P[319-:32]) - $signed(P[1357-:32])];
						FpRound = Mf[($signed(P[319-:32]) - $signed(P[1357-:32])) - 2];
					end
					2'h1: begin
						FpGuard = Mf[($signed(P[319-:32]) - $signed(P[1227-:32])) - 1];
						FpLsbRes = Mf[$signed(P[319-:32]) - $signed(P[1227-:32])];
						FpRound = Mf[($signed(P[319-:32]) - $signed(P[1227-:32])) - 2];
					end
					2'h0: begin
						FpGuard = Mf[($signed(P[319-:32]) - $signed(P[1097-:32])) - 1];
						FpLsbRes = Mf[$signed(P[319-:32]) - $signed(P[1097-:32])];
						FpRound = Mf[($signed(P[319-:32]) - $signed(P[1097-:32])) - 2];
					end
					2'h2: begin
						FpGuard = Mf[($signed(P[319-:32]) - $signed(P[967-:32])) - 1];
						FpLsbRes = Mf[$signed(P[319-:32]) - $signed(P[967-:32])];
						FpRound = Mf[($signed(P[319-:32]) - $signed(P[967-:32])) - 2];
					end
				endcase
			end
		end
	endgenerate
	assign Guard = (CvtToInt ? Mf[($signed(P[319-:32]) - $signed(P[4216-:32])) - 1] : FpGuard);
	assign LsbRes = (CvtToInt ? Mf[$signed(P[319-:32]) - $signed(P[4216-:32])] : FpLsbRes);
	assign Round = (CvtToInt ? Mf[($signed(P[319-:32]) - $signed(P[4216-:32])) - 2] : FpRound);
	always @(*) begin
		if (_sv2v_0)
			;
		case (Frm)
			3'b000: CalcPlus1 = Guard & ((Round | Sticky) | LsbRes);
			3'b001: CalcPlus1 = 1'b0;
			3'b010: CalcPlus1 = Ms;
			3'b011: CalcPlus1 = ~Ms;
			3'b100: CalcPlus1 = Guard;
			default: CalcPlus1 = 1'bx;
		endcase
		case (Frm)
			3'b000: UfCalcPlus1 = Round & (Sticky | Guard);
			3'b001: UfCalcPlus1 = 1'b0;
			3'b010: UfCalcPlus1 = Ms;
			3'b011: UfCalcPlus1 = ~Ms;
			3'b100: UfCalcPlus1 = Round;
			default: UfCalcPlus1 = 1'bx;
		endcase
	end
	assign Plus1 = CalcPlus1 & ((Sticky | Round) | Guard);
	assign FpPlus1 = Plus1 & ~CvtToInt;
	assign UfPlus1 = UfCalcPlus1 & (Sticky | Round);
	function automatic signed [(($signed(P[1389-:32]) + 1) + $signed(P[967-:32])) - 1:0] sv2v_cast_5E34A_signed;
		input reg signed [(($signed(P[1389-:32]) + 1) + $signed(P[967-:32])) - 1:0] inp;
		sv2v_cast_5E34A_signed = inp;
	endfunction
	function automatic signed [((($signed(P[1097-:32]) - $signed(P[967-:32])) - 2) >= 0 ? ($signed(P[1097-:32]) - $signed(P[967-:32])) - 1 : 3 - ($signed(P[1097-:32]) - $signed(P[967-:32]))) - 1:0] sv2v_cast_EF507_signed;
		input reg signed [((($signed(P[1097-:32]) - $signed(P[967-:32])) - 2) >= 0 ? ($signed(P[1097-:32]) - $signed(P[967-:32])) - 1 : 3 - ($signed(P[1097-:32]) - $signed(P[967-:32]))) - 1:0] inp;
		sv2v_cast_EF507_signed = inp;
	endfunction
	function automatic signed [((($signed(P[1227-:32]) - $signed(P[1097-:32])) - 2) >= 0 ? ($signed(P[1227-:32]) - $signed(P[1097-:32])) - 1 : 3 - ($signed(P[1227-:32]) - $signed(P[1097-:32]))) - 1:0] sv2v_cast_5435B_signed;
		input reg signed [((($signed(P[1227-:32]) - $signed(P[1097-:32])) - 2) >= 0 ? ($signed(P[1227-:32]) - $signed(P[1097-:32])) - 1 : 3 - ($signed(P[1227-:32]) - $signed(P[1097-:32]))) - 1:0] inp;
		sv2v_cast_5435B_signed = inp;
	endfunction
	function automatic signed [((($signed(P[1357-:32]) - $signed(P[1227-:32])) - 2) >= 0 ? ($signed(P[1357-:32]) - $signed(P[1227-:32])) - 1 : 3 - ($signed(P[1357-:32]) - $signed(P[1227-:32]))) - 1:0] sv2v_cast_8F6E9_signed;
		input reg signed [((($signed(P[1357-:32]) - $signed(P[1227-:32])) - 2) >= 0 ? ($signed(P[1357-:32]) - $signed(P[1227-:32])) - 1 : 3 - ($signed(P[1357-:32]) - $signed(P[1227-:32]))) - 1:0] inp;
		sv2v_cast_8F6E9_signed = inp;
	endfunction
	function automatic signed [(($signed(P[837-:32]) + 1) + $signed(P[481-:32])) - 1:0] sv2v_cast_34886_signed;
		input reg signed [(($signed(P[837-:32]) + 1) + $signed(P[481-:32])) - 1:0] inp;
		sv2v_cast_34886_signed = inp;
	endfunction
	function automatic signed [((($signed(P[611-:32]) - $signed(P[481-:32])) - 2) >= 0 ? ($signed(P[611-:32]) - $signed(P[481-:32])) - 1 : 3 - ($signed(P[611-:32]) - $signed(P[481-:32]))) - 1:0] sv2v_cast_3E459_signed;
		input reg signed [((($signed(P[611-:32]) - $signed(P[481-:32])) - 2) >= 0 ? ($signed(P[611-:32]) - $signed(P[481-:32])) - 1 : 3 - ($signed(P[611-:32]) - $signed(P[481-:32]))) - 1:0] inp;
		sv2v_cast_3E459_signed = inp;
	endfunction
	function automatic signed [((($signed(P[805-:32]) - $signed(P[611-:32])) - 2) >= 0 ? ($signed(P[805-:32]) - $signed(P[611-:32])) - 1 : 3 - ($signed(P[805-:32]) - $signed(P[611-:32]))) - 1:0] sv2v_cast_EB806_signed;
		input reg signed [((($signed(P[805-:32]) - $signed(P[611-:32])) - 2) >= 0 ? ($signed(P[805-:32]) - $signed(P[611-:32])) - 1 : 3 - ($signed(P[805-:32]) - $signed(P[611-:32]))) - 1:0] inp;
		sv2v_cast_EB806_signed = inp;
	endfunction
	function automatic signed [(($signed(P[837-:32]) + 1) + $signed(P[611-:32])) - 1:0] sv2v_cast_47E55_signed;
		input reg signed [(($signed(P[837-:32]) + 1) + $signed(P[611-:32])) - 1:0] inp;
		sv2v_cast_47E55_signed = inp;
	endfunction
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk3
			assign RoundAdd = {{$signed(P[901-:32]) {1'b0}}, FpPlus1};
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk3
			assign RoundAdd = {sv2v_cast_47E55_signed(0), FpPlus1 & ~OutFmt, sv2v_cast_EB806_signed(0), FpPlus1 & OutFmt};
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk3
			assign RoundAdd = {sv2v_cast_34886_signed(0), FpPlus1 & (OutFmt == P[449-:2]), sv2v_cast_3E459_signed(0), FpPlus1 & (OutFmt == P[579-:2]), sv2v_cast_EB806_signed(0), FpPlus1 & (OutFmt == P[773-:2])};
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk3
			assign RoundAdd = {sv2v_cast_5E34A_signed(0), FpPlus1 & (OutFmt == P[903-:2]), sv2v_cast_EF507_signed(0), FpPlus1 & (OutFmt == P[1033-:2]), sv2v_cast_5435B_signed(0), FpPlus1 & (OutFmt == P[1163-:2]), sv2v_cast_8F6E9_signed(0), FpPlus1 & (OutFmt == P[1293-:2])};
		end
	endgenerate
	assign RoundFrac = Mf[$signed(P[319-:32]) - 1:$signed(P[319-:32]) - $signed(P[805-:32])];
	always @(*) begin
		if (_sv2v_0)
			;
		case (PostProcSel)
			2'b10: Me = FmaMe;
			2'b00: Me = {CvtCe[$signed(P[837-:32])], CvtCe} & {$signed(P[837-:32]) + 2 {~CvtResSubnormUf | CvtResUf}};
			2'b01: Me = Ue;
			default: Me = 1'sb0;
		endcase
	end
	assign {FullRe, Rf} = {Me, RoundFrac} + RoundAdd;
	assign Re = FullRe[$signed(P[837-:32]) - 1:0];
	initial _sv2v_0 = 0;
endmodule
module roundsign (
	Xs,
	Ys,
	CvtCs,
	FmaSs,
	Sqrt,
	FmaOp,
	DivOp,
	CvtOp,
	Ms
);
	input wire Xs;
	input wire Ys;
	input wire CvtCs;
	input wire FmaSs;
	input wire Sqrt;
	input wire FmaOp;
	input wire DivOp;
	input wire CvtOp;
	output wire Ms;
	wire Qs;
	assign Qs = Xs ^ (Ys & ~Sqrt);
	assign Ms = ((FmaSs & FmaOp) | (CvtCs & CvtOp)) | (Qs & DivOp);
endmodule
module shiftcorrection (
	Shifted,
	DivOp,
	DivResSubnorm,
	DivUe,
	DivSubnormShiftPos,
	FmaOp,
	NormSumExp,
	FmaPreResultSubnorm,
	FmaSZero,
	FmaMe,
	Mf,
	Ue
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[319-:32]) - 1:0] Shifted;
	input wire DivOp;
	input wire DivResSubnorm;
	input wire [$signed(P[837-:32]) + 1:0] DivUe;
	input wire DivSubnormShiftPos;
	input wire FmaOp;
	input wire [$signed(P[837-:32]) + 1:0] NormSumExp;
	input wire FmaPreResultSubnorm;
	input wire FmaSZero;
	output wire [$signed(P[837-:32]) + 1:0] FmaMe;
	output reg [$signed(P[319-:32]) - 1:0] Mf;
	output wire [$signed(P[837-:32]) + 1:0] Ue;
	wire ResSubnorm;
	wire LZAPlus1;
	wire LeftShiftQm;
	wire RightShift;
	assign LZAPlus1 = Shifted[$signed(P[319-:32]) - 1];
	assign LeftShiftQm = LZAPlus1 | ((DivUe == 1) & ~LZAPlus1);
	assign RightShift = (FmaOp ? LZAPlus1 : LeftShiftQm);
	always @(*) begin
		if (_sv2v_0)
			;
		if (FmaOp | (DivOp & ~DivResSubnorm)) begin
			if (RightShift)
				Mf = {Shifted[$signed(P[319-:32]) - 2:1], 2'b00};
			else
				Mf = {Shifted[$signed(P[319-:32]) - 3:0], 2'b00};
		end
		else
			Mf = Shifted[$signed(P[319-:32]) - 1:0];
	end
	assign FmaMe = ((NormSumExp + {{$signed(P[837-:32]) + 1 {1'b0}}, LZAPlus1}) + {{$signed(P[837-:32]) + 1 {1'b0}}, FmaPreResultSubnorm}) & {$signed(P[837-:32]) + 2 {~(FmaSZero | ResSubnorm)}};
	assign ResSubnorm = (FmaPreResultSubnorm & ~Shifted[$signed(P[319-:32]) - 2]) & ~Shifted[$signed(P[319-:32]) - 1];
	function automatic signed [(($signed(P[837-:32]) + 0) >= 0 ? $signed(P[837-:32]) + 1 : 1 - ($signed(P[837-:32]) + 0)) - 1:0] sv2v_cast_97D7C_signed;
		input reg signed [(($signed(P[837-:32]) + 0) >= 0 ? $signed(P[837-:32]) + 1 : 1 - ($signed(P[837-:32]) + 0)) - 1:0] inp;
		sv2v_cast_97D7C_signed = inp;
	endfunction
	assign Ue = (DivResSubnorm & DivSubnormShiftPos ? 0 : DivUe - {sv2v_cast_97D7C_signed(0), ~LZAPlus1});
	initial _sv2v_0 = 0;
endmodule
module specialcase (
	Xs,
	Xm,
	Ym,
	Zm,
	XNaN,
	YNaN,
	ZNaN,
	Frm,
	OutFmt,
	InfIn,
	NaNIn,
	XInf,
	YInf,
	XZero,
	Plus1,
	Rs,
	Invalid,
	Overflow,
	Re,
	FullRe,
	Rf,
	FmaOp,
	DivOp,
	DivByZero,
	CvtOp,
	IntZero,
	IntToFp,
	Int64,
	Signed,
	Zfa,
	CvtCe,
	IntInvalid,
	CvtResUf,
	CvtNegRes,
	PostProcRes,
	FCvtIntRes
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire Xs;
	input wire [$signed(P[805-:32]):0] Xm;
	input wire [$signed(P[805-:32]):0] Ym;
	input wire [$signed(P[805-:32]):0] Zm;
	input wire XNaN;
	input wire YNaN;
	input wire ZNaN;
	input wire [2:0] Frm;
	input wire [$signed(P[707-:32]) - 1:0] OutFmt;
	input wire InfIn;
	input wire NaNIn;
	input wire XInf;
	input wire YInf;
	input wire XZero;
	input wire Plus1;
	input wire Rs;
	input wire Invalid;
	input wire Overflow;
	input wire [$signed(P[837-:32]) - 1:0] Re;
	input wire [$signed(P[837-:32]) + 1:0] FullRe;
	input wire [$signed(P[805-:32]) - 1:0] Rf;
	input wire FmaOp;
	input wire DivOp;
	input wire DivByZero;
	input wire CvtOp;
	input wire IntZero;
	input wire IntToFp;
	input wire Int64;
	input wire Signed;
	input wire Zfa;
	input wire [$signed(P[837-:32]):0] CvtCe;
	input wire IntInvalid;
	input wire CvtResUf;
	input wire [$signed(P[4216-:32]) + 1:0] CvtNegRes;
	output reg [$signed(P[901-:32]) - 1:0] PostProcRes;
	output reg [$signed(P[4216-:32]) - 1:0] FCvtIntRes;
	reg [$signed(P[901-:32]) - 1:0] XNaNRes;
	reg [$signed(P[901-:32]) - 1:0] YNaNRes;
	reg [$signed(P[901-:32]) - 1:0] ZNaNRes;
	reg [$signed(P[901-:32]) - 1:0] InvalidRes;
	reg [$signed(P[901-:32]) - 1:0] UfRes;
	reg [$signed(P[901-:32]) - 1:0] OfRes;
	reg [$signed(P[901-:32]) - 1:0] NormRes;
	reg [$signed(P[4216-:32]) - 1:0] OfIntRes;
	reg [$signed(P[4216-:32]) - 1:0] OfIntRes2;
	reg [$signed(P[4216-:32]) - 1:0] Int64Res;
	wire OfResMax;
	wire KillRes;
	wire SelOfRes;
	reg SelCvtOfRes;
	assign OfResMax = ((~InfIn | (IntToFp & CvtOp)) & ~DivByZero) & (((Frm[1:0] == 2'b01) | ((Frm[1:0] == 2'b10) & ~Rs)) | ((Frm[1:0] == 2'b11) & Rs));
	function automatic signed [(($signed(P[901-:32]) - 3) >= 0 ? $signed(P[901-:32]) - 2 : 4 - $signed(P[901-:32])) - 1:0] sv2v_cast_E1A99_signed;
		input reg signed [(($signed(P[901-:32]) - 3) >= 0 ? $signed(P[901-:32]) - 2 : 4 - $signed(P[901-:32])) - 1:0] inp;
		sv2v_cast_E1A99_signed = inp;
	endfunction
	function automatic signed [(($signed(P[1227-:32]) - 2) >= 0 ? $signed(P[1227-:32]) - 1 : 3 - $signed(P[1227-:32])) - 1:0] sv2v_cast_46E5E_signed;
		input reg signed [(($signed(P[1227-:32]) - 2) >= 0 ? $signed(P[1227-:32]) - 1 : 3 - $signed(P[1227-:32])) - 1:0] inp;
		sv2v_cast_46E5E_signed = inp;
	endfunction
	function automatic signed [$signed(P[1227-:32]) - 1:0] sv2v_cast_4FCCE_signed;
		input reg signed [$signed(P[1227-:32]) - 1:0] inp;
		sv2v_cast_4FCCE_signed = inp;
	endfunction
	function automatic signed [(($signed(P[1291-:32]) - 3) >= 0 ? $signed(P[1291-:32]) - 2 : 4 - $signed(P[1291-:32])) - 1:0] sv2v_cast_44A89_signed;
		input reg signed [(($signed(P[1291-:32]) - 3) >= 0 ? $signed(P[1291-:32]) - 2 : 4 - $signed(P[1291-:32])) - 1:0] inp;
		sv2v_cast_44A89_signed = inp;
	endfunction
	function automatic signed [(($signed(P[1097-:32]) - 2) >= 0 ? $signed(P[1097-:32]) - 1 : 3 - $signed(P[1097-:32])) - 1:0] sv2v_cast_B8EE9_signed;
		input reg signed [(($signed(P[1097-:32]) - 2) >= 0 ? $signed(P[1097-:32]) - 1 : 3 - $signed(P[1097-:32])) - 1:0] inp;
		sv2v_cast_B8EE9_signed = inp;
	endfunction
	function automatic signed [$signed(P[1097-:32]) - 1:0] sv2v_cast_CACF9_signed;
		input reg signed [$signed(P[1097-:32]) - 1:0] inp;
		sv2v_cast_CACF9_signed = inp;
	endfunction
	function automatic signed [(($signed(P[1161-:32]) - 3) >= 0 ? $signed(P[1161-:32]) - 2 : 4 - $signed(P[1161-:32])) - 1:0] sv2v_cast_C389E_signed;
		input reg signed [(($signed(P[1161-:32]) - 3) >= 0 ? $signed(P[1161-:32]) - 2 : 4 - $signed(P[1161-:32])) - 1:0] inp;
		sv2v_cast_C389E_signed = inp;
	endfunction
	function automatic signed [(($signed(P[967-:32]) - 2) >= 0 ? $signed(P[967-:32]) - 1 : 3 - $signed(P[967-:32])) - 1:0] sv2v_cast_67652_signed;
		input reg signed [(($signed(P[967-:32]) - 2) >= 0 ? $signed(P[967-:32]) - 1 : 3 - $signed(P[967-:32])) - 1:0] inp;
		sv2v_cast_67652_signed = inp;
	endfunction
	function automatic signed [$signed(P[967-:32]) - 1:0] sv2v_cast_17AC2_signed;
		input reg signed [$signed(P[967-:32]) - 1:0] inp;
		sv2v_cast_17AC2_signed = inp;
	endfunction
	function automatic signed [(($signed(P[1031-:32]) - 3) >= 0 ? $signed(P[1031-:32]) - 2 : 4 - $signed(P[1031-:32])) - 1:0] sv2v_cast_E3205_signed;
		input reg signed [(($signed(P[1031-:32]) - 3) >= 0 ? $signed(P[1031-:32]) - 2 : 4 - $signed(P[1031-:32])) - 1:0] inp;
		sv2v_cast_E3205_signed = inp;
	endfunction
	function automatic signed [(($signed(P[611-:32]) - 2) >= 0 ? $signed(P[611-:32]) - 1 : 3 - $signed(P[611-:32])) - 1:0] sv2v_cast_B7E13_signed;
		input reg signed [(($signed(P[611-:32]) - 2) >= 0 ? $signed(P[611-:32]) - 1 : 3 - $signed(P[611-:32])) - 1:0] inp;
		sv2v_cast_B7E13_signed = inp;
	endfunction
	function automatic signed [$signed(P[611-:32]) - 1:0] sv2v_cast_C55D7_signed;
		input reg signed [$signed(P[611-:32]) - 1:0] inp;
		sv2v_cast_C55D7_signed = inp;
	endfunction
	function automatic signed [(($signed(P[675-:32]) - 3) >= 0 ? $signed(P[675-:32]) - 2 : 4 - $signed(P[675-:32])) - 1:0] sv2v_cast_4EE8E_signed;
		input reg signed [(($signed(P[675-:32]) - 3) >= 0 ? $signed(P[675-:32]) - 2 : 4 - $signed(P[675-:32])) - 1:0] inp;
		sv2v_cast_4EE8E_signed = inp;
	endfunction
	function automatic signed [(($signed(P[481-:32]) - 2) >= 0 ? $signed(P[481-:32]) - 1 : 3 - $signed(P[481-:32])) - 1:0] sv2v_cast_E1570_signed;
		input reg signed [(($signed(P[481-:32]) - 2) >= 0 ? $signed(P[481-:32]) - 1 : 3 - $signed(P[481-:32])) - 1:0] inp;
		sv2v_cast_E1570_signed = inp;
	endfunction
	function automatic signed [$signed(P[481-:32]) - 1:0] sv2v_cast_69944_signed;
		input reg signed [$signed(P[481-:32]) - 1:0] inp;
		sv2v_cast_69944_signed = inp;
	endfunction
	function automatic signed [(($signed(P[545-:32]) - 3) >= 0 ? $signed(P[545-:32]) - 2 : 4 - $signed(P[545-:32])) - 1:0] sv2v_cast_2D6DD_signed;
		input reg signed [(($signed(P[545-:32]) - 3) >= 0 ? $signed(P[545-:32]) - 2 : 4 - $signed(P[545-:32])) - 1:0] inp;
		sv2v_cast_2D6DD_signed = inp;
	endfunction
	function automatic signed [$signed(P[901-:32]) - 1:0] sv2v_cast_7604C_signed;
		input reg signed [$signed(P[901-:32]) - 1:0] inp;
		sv2v_cast_7604C_signed = inp;
	endfunction
	generate
		if ($signed(P[739-:32]) == 1) begin : genblk1
			if (P[4184]) begin : genblk1
				wire [$signed(P[901-:32]):1] sv2v_tmp_0825B;
				assign sv2v_tmp_0825B = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:0]};
				always @(*) XNaNRes = sv2v_tmp_0825B;
				wire [$signed(P[901-:32]):1] sv2v_tmp_3B8DB;
				assign sv2v_tmp_3B8DB = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, Ym[$signed(P[805-:32]) - 2:0]};
				always @(*) YNaNRes = sv2v_tmp_3B8DB;
				wire [$signed(P[901-:32]):1] sv2v_tmp_6789B;
				assign sv2v_tmp_6789B = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, Zm[$signed(P[805-:32]) - 2:0]};
				always @(*) ZNaNRes = sv2v_tmp_6789B;
				wire [$signed(P[901-:32]):1] sv2v_tmp_4F543;
				assign sv2v_tmp_4F543 = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, {$signed(P[805-:32]) - 1 {1'b0}}};
				always @(*) InvalidRes = sv2v_tmp_4F543;
			end
			else begin : genblk1
				wire [$signed(P[901-:32]):1] sv2v_tmp_4F543;
				assign sv2v_tmp_4F543 = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, {$signed(P[805-:32]) - 1 {1'b0}}};
				always @(*) InvalidRes = sv2v_tmp_4F543;
			end
			wire [$signed(P[901-:32]):1] sv2v_tmp_9A5CB;
			assign sv2v_tmp_9A5CB = (OfResMax ? {Rs, {$signed(P[837-:32]) - 1 {1'b1}}, 1'b0, {$signed(P[805-:32]) {1'b1}}} : {Rs, {$signed(P[837-:32]) {1'b1}}, {$signed(P[805-:32]) {1'b0}}});
			always @(*) OfRes = sv2v_tmp_9A5CB;
			wire [$signed(P[901-:32]):1] sv2v_tmp_33538;
			assign sv2v_tmp_33538 = {Rs, {$signed(P[901-:32]) - 2 {1'b0}}, (Plus1 & Frm[1]) & ~(DivOp & YInf)};
			always @(*) UfRes = sv2v_tmp_33538;
			wire [$signed(P[901-:32]):1] sv2v_tmp_3EE80;
			assign sv2v_tmp_3EE80 = {Rs, Re, Rf};
			always @(*) NormRes = sv2v_tmp_3EE80;
		end
		else if ($signed(P[739-:32]) == 2) begin : genblk1
			if (P[4184]) begin : genblk1
				wire [$signed(P[901-:32]):1] sv2v_tmp_69DFA;
				assign sv2v_tmp_69DFA = (OutFmt ? {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:0]} : {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 1'b0, {$signed(P[643-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[611-:32])]});
				always @(*) XNaNRes = sv2v_tmp_69DFA;
				wire [$signed(P[901-:32]):1] sv2v_tmp_9717B;
				assign sv2v_tmp_9717B = (OutFmt ? {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, Ym[$signed(P[805-:32]) - 2:0]} : {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 1'b0, {$signed(P[643-:32]) {1'b1}}, 1'b1, Ym[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[611-:32])]});
				always @(*) YNaNRes = sv2v_tmp_9717B;
				wire [$signed(P[901-:32]):1] sv2v_tmp_19F38;
				assign sv2v_tmp_19F38 = (OutFmt ? {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, Zm[$signed(P[805-:32]) - 2:0]} : {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 1'b0, {$signed(P[643-:32]) {1'b1}}, 1'b1, Zm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[611-:32])]});
				always @(*) ZNaNRes = sv2v_tmp_19F38;
				wire [$signed(P[901-:32]):1] sv2v_tmp_5B3B4;
				assign sv2v_tmp_5B3B4 = (OutFmt ? {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, {$signed(P[805-:32]) - 1 {1'b0}}} : {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 1'b0, {$signed(P[643-:32]) {1'b1}}, 1'b1, sv2v_cast_B7E13_signed(0)});
				always @(*) InvalidRes = sv2v_tmp_5B3B4;
			end
			else begin : genblk1
				wire [$signed(P[901-:32]):1] sv2v_tmp_5B3B4;
				assign sv2v_tmp_5B3B4 = (OutFmt ? {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, {$signed(P[805-:32]) - 1 {1'b0}}} : {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 1'b0, {$signed(P[643-:32]) {1'b1}}, 1'b1, sv2v_cast_B7E13_signed(0)});
				always @(*) InvalidRes = sv2v_tmp_5B3B4;
			end
			always @(*) begin
				if (_sv2v_0)
					;
				if (OutFmt) begin
					if (OfResMax)
						OfRes = {Rs, {$signed(P[837-:32]) - 1 {1'b1}}, 1'b0, {$signed(P[805-:32]) {1'b1}}};
					else
						OfRes = {Rs, {$signed(P[837-:32]) {1'b1}}, {$signed(P[805-:32]) {1'b0}}};
				end
				else if (OfResMax)
					OfRes = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, Rs, {$signed(P[643-:32]) - 1 {1'b1}}, 1'b0, {$signed(P[611-:32]) {1'b1}}};
				else
					OfRes = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, Rs, {$signed(P[643-:32]) {1'b1}}, sv2v_cast_C55D7_signed(0)};
			end
			wire [$signed(P[901-:32]):1] sv2v_tmp_E2FF3;
			assign sv2v_tmp_E2FF3 = (OutFmt ? {Rs, sv2v_cast_E1A99_signed(0), (Plus1 & Frm[1]) & ~(DivOp & YInf)} : {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, Rs, sv2v_cast_4EE8E_signed(0), (Plus1 & Frm[1]) & ~(DivOp & YInf)});
			always @(*) UfRes = sv2v_tmp_E2FF3;
			wire [$signed(P[901-:32]):1] sv2v_tmp_682A4;
			assign sv2v_tmp_682A4 = (OutFmt ? {Rs, Re, Rf} : {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, Rs, Re[$signed(P[643-:32]) - 1:0], Rf[$signed(P[805-:32]) - 1:$signed(P[805-:32]) - $signed(P[611-:32])]});
			always @(*) NormRes = sv2v_tmp_682A4;
		end
		else if ($signed(P[739-:32]) == 3) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				case (OutFmt)
					P[773-:2]: begin
						if (P[4184]) begin
							XNaNRes = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:0]};
							YNaNRes = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, Ym[$signed(P[805-:32]) - 2:0]};
							ZNaNRes = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, Zm[$signed(P[805-:32]) - 2:0]};
							InvalidRes = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, {$signed(P[805-:32]) - 1 {1'b0}}};
						end
						else
							InvalidRes = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, {$signed(P[805-:32]) - 1 {1'b0}}};
						OfRes = (OfResMax ? {Rs, {$signed(P[837-:32]) - 1 {1'b1}}, 1'b0, {$signed(P[805-:32]) {1'b1}}} : {Rs, {$signed(P[837-:32]) {1'b1}}, {$signed(P[805-:32]) {1'b0}}});
						UfRes = {Rs, sv2v_cast_E1A99_signed(0), (Plus1 & Frm[1]) & ~(DivOp & YInf)};
						NormRes = {Rs, Re, Rf};
					end
					P[579-:2]: begin
						if (P[4184]) begin
							XNaNRes = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 1'b0, {$signed(P[643-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[611-:32])]};
							YNaNRes = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 1'b0, {$signed(P[643-:32]) {1'b1}}, 1'b1, Ym[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[611-:32])]};
							ZNaNRes = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 1'b0, {$signed(P[643-:32]) {1'b1}}, 1'b1, Zm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[611-:32])]};
							InvalidRes = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 1'b0, {$signed(P[643-:32]) {1'b1}}, 1'b1, sv2v_cast_B7E13_signed(0)};
						end
						else
							InvalidRes = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, 1'b0, {$signed(P[643-:32]) {1'b1}}, 1'b1, sv2v_cast_B7E13_signed(0)};
						OfRes = (OfResMax ? {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, Rs, {$signed(P[643-:32]) - 1 {1'b1}}, 1'b0, {$signed(P[611-:32]) {1'b1}}} : {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, Rs, {$signed(P[643-:32]) {1'b1}}, sv2v_cast_C55D7_signed(0)});
						UfRes = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, Rs, sv2v_cast_4EE8E_signed(0), (Plus1 & Frm[1]) & ~(DivOp & YInf)};
						NormRes = {{$signed(P[901-:32]) - $signed(P[675-:32]) {1'b1}}, Rs, Re[$signed(P[643-:32]) - 1:0], Rf[$signed(P[805-:32]) - 1:$signed(P[805-:32]) - $signed(P[611-:32])]};
					end
					P[449-:2]: begin
						if (P[4184]) begin
							XNaNRes = {{$signed(P[901-:32]) - $signed(P[545-:32]) {1'b1}}, 1'b0, {$signed(P[513-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[481-:32])]};
							YNaNRes = {{$signed(P[901-:32]) - $signed(P[545-:32]) {1'b1}}, 1'b0, {$signed(P[513-:32]) {1'b1}}, 1'b1, Ym[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[481-:32])]};
							ZNaNRes = {{$signed(P[901-:32]) - $signed(P[545-:32]) {1'b1}}, 1'b0, {$signed(P[513-:32]) {1'b1}}, 1'b1, Zm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[481-:32])]};
							InvalidRes = {{$signed(P[901-:32]) - $signed(P[545-:32]) {1'b1}}, 1'b0, {$signed(P[513-:32]) {1'b1}}, 1'b1, sv2v_cast_E1570_signed(0)};
						end
						else
							InvalidRes = {{$signed(P[901-:32]) - $signed(P[545-:32]) {1'b1}}, 1'b0, {$signed(P[513-:32]) {1'b1}}, 1'b1, sv2v_cast_E1570_signed(0)};
						OfRes = (OfResMax ? {{$signed(P[901-:32]) - $signed(P[545-:32]) {1'b1}}, Rs, {$signed(P[513-:32]) - 1 {1'b1}}, 1'b0, {$signed(P[481-:32]) {1'b1}}} : {{$signed(P[901-:32]) - $signed(P[545-:32]) {1'b1}}, Rs, {$signed(P[513-:32]) {1'b1}}, sv2v_cast_69944_signed(0)});
						UfRes = {{$signed(P[901-:32]) - $signed(P[545-:32]) {1'b1}}, Rs, sv2v_cast_2D6DD_signed(0), (Plus1 & Frm[1]) & ~(DivOp & YInf)};
						NormRes = {{$signed(P[901-:32]) - $signed(P[545-:32]) {1'b1}}, Rs, Re[$signed(P[513-:32]) - 1:0], Rf[$signed(P[805-:32]) - 1:$signed(P[805-:32]) - $signed(P[481-:32])]};
					end
					default: begin
						if (P[4184]) begin
							XNaNRes = sv2v_cast_7604C_signed(0);
							YNaNRes = sv2v_cast_7604C_signed(0);
							ZNaNRes = sv2v_cast_7604C_signed(0);
							InvalidRes = sv2v_cast_7604C_signed(0);
						end
						else
							InvalidRes = sv2v_cast_7604C_signed(0);
						OfRes = sv2v_cast_7604C_signed(0);
						UfRes = sv2v_cast_7604C_signed(0);
						NormRes = sv2v_cast_7604C_signed(0);
					end
				endcase
			end
		end
		else if ($signed(P[739-:32]) == 4) begin : genblk1
			always @(*) begin
				if (_sv2v_0)
					;
				case (OutFmt)
					2'h3: begin
						if (P[4184]) begin
							XNaNRes = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:0]};
							YNaNRes = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, Ym[$signed(P[805-:32]) - 2:0]};
							ZNaNRes = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, Zm[$signed(P[805-:32]) - 2:0]};
							InvalidRes = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, {$signed(P[805-:32]) - 1 {1'b0}}};
						end
						else
							InvalidRes = {1'b0, {$signed(P[837-:32]) {1'b1}}, 1'b1, {$signed(P[805-:32]) - 1 {1'b0}}};
						OfRes = (OfResMax ? {Rs, {$signed(P[837-:32]) - 1 {1'b1}}, 1'b0, {$signed(P[805-:32]) {1'b1}}} : {Rs, {$signed(P[837-:32]) {1'b1}}, {$signed(P[805-:32]) {1'b0}}});
						UfRes = {Rs, sv2v_cast_E1A99_signed(0), (Plus1 & Frm[1]) & ~(DivOp & YInf)};
						NormRes = {Rs, Re, Rf};
					end
					2'h1: begin
						if (P[4184]) begin
							XNaNRes = {{$signed(P[901-:32]) - $signed(P[1291-:32]) {1'b1}}, 1'b0, {$signed(P[1259-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[1227-:32])]};
							YNaNRes = {{$signed(P[901-:32]) - $signed(P[1291-:32]) {1'b1}}, 1'b0, {$signed(P[1259-:32]) {1'b1}}, 1'b1, Ym[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[1227-:32])]};
							ZNaNRes = {{$signed(P[901-:32]) - $signed(P[1291-:32]) {1'b1}}, 1'b0, {$signed(P[1259-:32]) {1'b1}}, 1'b1, Zm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[1227-:32])]};
							InvalidRes = {{$signed(P[901-:32]) - $signed(P[1291-:32]) {1'b1}}, 1'b0, {$signed(P[1259-:32]) {1'b1}}, 1'b1, sv2v_cast_46E5E_signed(0)};
						end
						else
							InvalidRes = {{$signed(P[901-:32]) - $signed(P[1291-:32]) {1'b1}}, 1'b0, {$signed(P[1259-:32]) {1'b1}}, 1'b1, sv2v_cast_46E5E_signed(0)};
						OfRes = (OfResMax ? {{$signed(P[901-:32]) - $signed(P[1291-:32]) {1'b1}}, Rs, {$signed(P[1259-:32]) - 1 {1'b1}}, 1'b0, {$signed(P[1227-:32]) {1'b1}}} : {{$signed(P[901-:32]) - $signed(P[1291-:32]) {1'b1}}, Rs, {$signed(P[1259-:32]) {1'b1}}, sv2v_cast_4FCCE_signed(0)});
						UfRes = {{$signed(P[901-:32]) - $signed(P[1291-:32]) {1'b1}}, Rs, sv2v_cast_44A89_signed(0), (Plus1 & Frm[1]) & ~(DivOp & YInf)};
						NormRes = {{$signed(P[901-:32]) - $signed(P[1291-:32]) {1'b1}}, Rs, Re[$signed(P[1259-:32]) - 1:0], Rf[$signed(P[805-:32]) - 1:$signed(P[805-:32]) - $signed(P[1227-:32])]};
					end
					2'h0: begin
						if (P[4184]) begin
							XNaNRes = {{$signed(P[901-:32]) - $signed(P[1161-:32]) {1'b1}}, 1'b0, {$signed(P[1129-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[1097-:32])]};
							YNaNRes = {{$signed(P[901-:32]) - $signed(P[1161-:32]) {1'b1}}, 1'b0, {$signed(P[1129-:32]) {1'b1}}, 1'b1, Ym[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[1097-:32])]};
							ZNaNRes = {{$signed(P[901-:32]) - $signed(P[1161-:32]) {1'b1}}, 1'b0, {$signed(P[1129-:32]) {1'b1}}, 1'b1, Zm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[1097-:32])]};
							InvalidRes = {{$signed(P[901-:32]) - $signed(P[1161-:32]) {1'b1}}, 1'b0, {$signed(P[1129-:32]) {1'b1}}, 1'b1, sv2v_cast_B8EE9_signed(0)};
						end
						else
							InvalidRes = {{$signed(P[901-:32]) - $signed(P[1161-:32]) {1'b1}}, 1'b0, {$signed(P[1129-:32]) {1'b1}}, 1'b1, sv2v_cast_B8EE9_signed(0)};
						OfRes = (OfResMax ? {{$signed(P[901-:32]) - $signed(P[1161-:32]) {1'b1}}, Rs, {$signed(P[1129-:32]) - 1 {1'b1}}, 1'b0, {$signed(P[1097-:32]) {1'b1}}} : {{$signed(P[901-:32]) - $signed(P[1161-:32]) {1'b1}}, Rs, {$signed(P[1129-:32]) {1'b1}}, sv2v_cast_CACF9_signed(0)});
						UfRes = {{$signed(P[901-:32]) - $signed(P[1161-:32]) {1'b1}}, Rs, sv2v_cast_C389E_signed(0), (Plus1 & Frm[1]) & ~(DivOp & YInf)};
						NormRes = {{$signed(P[901-:32]) - $signed(P[1161-:32]) {1'b1}}, Rs, Re[$signed(P[1129-:32]) - 1:0], Rf[$signed(P[805-:32]) - 1:$signed(P[805-:32]) - $signed(P[1097-:32])]};
					end
					2'h2: begin
						if (P[4184]) begin
							XNaNRes = {{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, 1'b0, {$signed(P[999-:32]) {1'b1}}, 1'b1, Xm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[967-:32])]};
							YNaNRes = {{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, 1'b0, {$signed(P[999-:32]) {1'b1}}, 1'b1, Ym[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[967-:32])]};
							ZNaNRes = {{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, 1'b0, {$signed(P[999-:32]) {1'b1}}, 1'b1, Zm[$signed(P[805-:32]) - 2:$signed(P[805-:32]) - $signed(P[967-:32])]};
							InvalidRes = {{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, 1'b0, {$signed(P[999-:32]) {1'b1}}, 1'b1, sv2v_cast_67652_signed(0)};
						end
						else
							InvalidRes = {{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, 1'b0, {$signed(P[999-:32]) {1'b1}}, 1'b1, sv2v_cast_67652_signed(0)};
						OfRes = (OfResMax ? {{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, Rs, {$signed(P[999-:32]) - 1 {1'b1}}, 1'b0, {$signed(P[967-:32]) {1'b1}}} : {{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, Rs, {$signed(P[999-:32]) {1'b1}}, sv2v_cast_17AC2_signed(0)});
						UfRes = {{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, Rs, sv2v_cast_E3205_signed(0), (Plus1 & Frm[1]) & ~(DivOp & YInf)};
						NormRes = {{$signed(P[901-:32]) - $signed(P[1031-:32]) {1'b1}}, Rs, Re[$signed(P[999-:32]) - 1:0], Rf[$signed(P[805-:32]) - 1:$signed(P[805-:32]) - $signed(P[967-:32])]};
					end
				endcase
			end
		end
	endgenerate
	assign KillRes = (CvtOp ? (CvtResUf | (XZero & ~IntToFp)) | (IntZero & IntToFp) : FullRe[$signed(P[837-:32]) + 1] | (((YInf & ~XInf) | XZero) & DivOp));
	assign SelOfRes = (Overflow | DivByZero) | (InfIn & ~(YInf & DivOp));
	generate
		if (P[4184]) begin : genblk2
			always @(*) begin
				if (_sv2v_0)
					;
				if (XNaN & ~(IntToFp & CvtOp))
					PostProcRes = XNaNRes;
				else if (YNaN & ~CvtOp)
					PostProcRes = YNaNRes;
				else if (ZNaN & FmaOp)
					PostProcRes = ZNaNRes;
				else if (Invalid)
					PostProcRes = InvalidRes;
				else if (SelOfRes)
					PostProcRes = OfRes;
				else if (KillRes)
					PostProcRes = UfRes;
				else
					PostProcRes = NormRes;
			end
		end
		else begin : genblk2
			always @(*) begin
				if (_sv2v_0)
					;
				if (NaNIn | Invalid)
					PostProcRes = InvalidRes;
				else if (SelOfRes)
					PostProcRes = OfRes;
				else if (KillRes)
					PostProcRes = UfRes;
				else
					PostProcRes = NormRes;
			end
		end
		if (P[4184]) begin : genblk3
			always @(*) begin
				if (_sv2v_0)
					;
				if (Signed) begin
					if (Xs & ~NaNIn) begin
						if (Int64)
							OfIntRes = {1'b1, {$signed(P[4216-:32]) - 1 {1'b0}}};
						else
							OfIntRes = {{$signed(P[4216-:32]) - 32 {1'b1}}, 1'b1, {31 {1'b0}}};
					end
					else if (Int64)
						OfIntRes = {1'b1, {$signed(P[4216-:32]) - 1 {1'b0}}};
					else
						OfIntRes = {{$signed(P[4216-:32]) - 32 {1'b1}}, 1'b1, {31 {1'b0}}};
				end
				else if (Xs & ~NaNIn)
					OfIntRes = {$signed(P[4216-:32]) {1'b1}};
				else
					OfIntRes = {$signed(P[4216-:32]) {1'b1}};
			end
		end
		else begin : genblk3
			always @(*) begin
				if (_sv2v_0)
					;
				if (Signed) begin
					if (Xs & ~NaNIn) begin
						if (Int64)
							OfIntRes = {1'b1, {$signed(P[4216-:32]) - 1 {1'b0}}};
						else
							OfIntRes = {{$signed(P[4216-:32]) - 32 {1'b1}}, 1'b1, {31 {1'b0}}};
					end
					else if (Int64)
						OfIntRes = {1'b0, {$signed(P[4216-:32]) - 1 {1'b1}}};
					else
						OfIntRes = {{$signed(P[4216-:32]) - 32 {1'b0}}, 1'b0, {31 {1'b1}}};
				end
				else if (Xs & ~NaNIn)
					OfIntRes = {$signed(P[4216-:32]) {1'b0}};
				else
					OfIntRes = {$signed(P[4216-:32]) {1'b1}};
			end
		end
		if (P[4069] & P[1493]) begin : genblk4
			always @(*) begin
				if (_sv2v_0)
					;
				if (Zfa)
					OfIntRes2 = 1'sb0;
				else
					OfIntRes2 = OfIntRes;
				if (Zfa)
					Int64Res = {{$signed(P[4216-:32]) - 32 {CvtNegRes[$signed(P[4216-:32]) - 1]}}, CvtNegRes[31:0]};
				else
					Int64Res = CvtNegRes[$signed(P[4216-:32]) - 1:0];
				if (Zfa)
					SelCvtOfRes = (InfIn | NaNIn) | (CvtCe > 84);
				else
					SelCvtOfRes = IntInvalid;
			end
		end
		else begin : genblk4
			always @(*) begin
				if (_sv2v_0)
					;
				OfIntRes2 = OfIntRes;
				Int64Res = CvtNegRes[$signed(P[4216-:32]) - 1:0];
				SelCvtOfRes = IntInvalid;
			end
		end
	endgenerate
	always @(*) begin
		if (_sv2v_0)
			;
		if (SelCvtOfRes)
			FCvtIntRes = OfIntRes2;
		else if (CvtCe[$signed(P[837-:32])]) begin
			if ((Xs & Signed) & Plus1)
				FCvtIntRes = {$signed(P[4216-:32]) {1'b1}};
			else
				FCvtIntRes = {{$signed(P[4216-:32]) - 1 {1'b0}}, Plus1};
		end
		else if (Int64)
			FCvtIntRes = Int64Res;
		else
			FCvtIntRes = {{$signed(P[4216-:32]) - 32 {CvtNegRes[31]}}, CvtNegRes[31:0]};
	end
	initial _sv2v_0 = 0;
endmodule
module flop (
	clk,
	d,
	q
);
	parameter WIDTH = 8;
	input wire clk;
	input wire [WIDTH - 1:0] d;
	output reg [WIDTH - 1:0] q;
	always @(posedge clk) q <= d;
endmodule
module flopen (
	clk,
	en,
	d,
	q
);
	parameter WIDTH = 8;
	input wire clk;
	input wire en;
	input wire [WIDTH - 1:0] d;
	output reg [WIDTH - 1:0] q;
	always @(posedge clk)
		if (en)
			q <= d;
endmodule
module flopenl (
	clk,
	load,
	en,
	d,
	val,
	q
);
	parameter WIDTH = 8;
	input wire clk;
	input wire load;
	input wire en;
	input wire [WIDTH - 1:0] d;
	input wire [WIDTH - 1:0] val;
	output reg [WIDTH - 1:0] q;
	always @(posedge clk)
		if (load)
			q <= val;
		else if (en)
			q <= d;
endmodule
module flopenl_8C148 (
	clk,
	load,
	en,
	d,
	val,
	q
);
	parameter WIDTH = 8;
	input wire clk;
	input wire load;
	input wire en;
	input wire [1:0] d;
	input wire [1:0] val;
	output reg [1:0] q;
	always @(posedge clk)
		if (load)
			q <= val;
		else if (en)
			q <= d;
endmodule
module flopenl_FC78A (
	clk,
	load,
	en,
	d,
	val,
	q
);
	parameter WIDTH = 8;
	input wire clk;
	input wire load;
	input wire en;
	input wire [3:0] d;
	input wire [3:0] val;
	output reg [3:0] q;
	always @(posedge clk)
		if (load)
			q <= val;
		else if (en)
			q <= d;
endmodule
module flopenr (
	clk,
	reset,
	en,
	d,
	q
);
	parameter WIDTH = 8;
	input wire clk;
	input wire reset;
	input wire en;
	input wire [WIDTH - 1:0] d;
	output reg [WIDTH - 1:0] q;
	always @(posedge clk)
		if (reset)
			q <= 1'sb0;
		else if (en)
			q <= d;
endmodule
module flopenrc (
	clk,
	reset,
	clear,
	en,
	d,
	q
);
	parameter WIDTH = 8;
	input wire clk;
	input wire reset;
	input wire clear;
	input wire en;
	input wire [WIDTH - 1:0] d;
	output reg [WIDTH - 1:0] q;
	always @(posedge clk)
		if (reset)
			q <= 1'sb0;
		else if (en) begin
			if (clear)
				q <= 1'sb0;
			else
				q <= d;
		end
endmodule
module flopr (
	clk,
	reset,
	d,
	q
);
	parameter WIDTH = 8;
	input wire clk;
	input wire reset;
	input wire [WIDTH - 1:0] d;
	output reg [WIDTH - 1:0] q;
	always @(posedge clk)
		if (reset)
			q <= 1'sb0;
		else
			q <= d;
endmodule
module synchronizer (
	clk,
	d,
	q
);
	input wire clk;
	input wire d;
	output reg q;
	reg mid;
	always @(posedge clk) begin
		mid <= d;
		q <= mid;
	end
endmodule
module ram1p1rwbe (
	clk,
	ce,
	addr,
	din,
	we,
	bwe,
	dout
);
	parameter USE_SRAM = 0;
	parameter DEPTH = 64;
	parameter WIDTH = 44;
	parameter PRELOAD_ENABLED = 0;
	input wire clk;
	input wire ce;
	input wire [$clog2(DEPTH) - 1:0] addr;
	input wire [WIDTH - 1:0] din;
	input wire we;
	input wire [(WIDTH - 1) / 8:0] bwe;
	output wire [WIDTH - 1:0] dout;
	generate
		if (((USE_SRAM == 1) & (WIDTH == 128)) & (DEPTH == 64)) begin : genblk1
			genvar _gv_index_8;
			wire [WIDTH - 1:0] BitWriteMask;
			for (_gv_index_8 = 0; _gv_index_8 < WIDTH; _gv_index_8 = _gv_index_8 + 1) begin : genblk1
				localparam index = _gv_index_8;
				assign BitWriteMask[index] = bwe[index / 8];
			end
			ram1p1rwbe_64x128 sram1A(
				.CLK(clk),
				.CEB(~ce),
				.WEB(~we),
				.A(addr),
				.D(din),
				.BWEB(~BitWriteMask),
				.Q(dout)
			);
		end
		else if (((USE_SRAM == 1) & (WIDTH == 44)) & (DEPTH == 64)) begin : genblk1
			genvar _gv_index_9;
			wire [WIDTH - 1:0] BitWriteMask;
			for (_gv_index_9 = 0; _gv_index_9 < WIDTH; _gv_index_9 = _gv_index_9 + 1) begin : genblk1
				localparam index = _gv_index_9;
				assign BitWriteMask[index] = bwe[index / 8];
			end
			ram1p1rwbe_64x44 sram1B(
				.CLK(clk),
				.CEB(~ce),
				.WEB(~we),
				.A(addr),
				.D(din),
				.BWEB(~BitWriteMask),
				.Q(dout)
			);
		end
		else if (((USE_SRAM == 1) & (WIDTH == 22)) & (DEPTH == 64)) begin : genblk1
			genvar _gv_index_10;
			wire [WIDTH - 1:0] BitWriteMask;
			for (_gv_index_10 = 0; _gv_index_10 < WIDTH; _gv_index_10 = _gv_index_10 + 1) begin : genblk1
				localparam index = _gv_index_10;
				assign BitWriteMask[index] = bwe[index / 8];
			end
			ram1p1rwbe_64x22 sram1B(
				.CLK(clk),
				.CEB(~ce),
				.WEB(~we),
				.A(addr),
				.D(din),
				.BWEB(~BitWriteMask),
				.Q(dout)
			);
		end
		else begin : ram
			reg [WIDTH - 1:0] RAM [DEPTH - 1:0];
			initial if (PRELOAD_ENABLED) begin
				if (WIDTH == 64)
					$readmemh({"$WALLY/fpga/src/data.mem"}, RAM, 0);
				else
					RAM[0] = 'h2197;
			end
			wire [$clog2(DEPTH) - 1:0] addrd;
			flopen #(.WIDTH($clog2(DEPTH))) adrreg(
				.clk(clk),
				.en(ce),
				.d(addr),
				.q(addrd)
			);
			assign dout = RAM[addrd];
			if (WIDTH >= 8) begin : genblk1
				integer i;
				always @(posedge clk)
					if (ce & we) begin
						for (i = 0; i < (WIDTH / 8); i = i + 1)
							if (bwe[i])
								RAM[addr][i * 8+:8] <= din[i * 8+:8];
					end
			end
			if ((WIDTH % 8) != 0) begin : genblk2
				always @(posedge clk)
					if ((ce & we) & bwe[WIDTH / 8])
						RAM[addr][WIDTH - 1:WIDTH - (WIDTH % 8)] <= din[WIDTH - 1:WIDTH - (WIDTH % 8)];
			end
		end
	endgenerate
endmodule
module ram1p1rwbe_64x128 (
	CLK,
	CEB,
	WEB,
	A,
	D,
	BWEB,
	Q
);
	input wire CLK;
	input wire CEB;
	input wire WEB;
	input wire [5:0] A;
	input wire [127:0] D;
	input wire [127:0] BWEB;
	output wire [127:0] Q;
	TS1N28HPCPSVTB64X128M4SW sramIP(
		.CLK(CLK),
		.CEB(CEB),
		.WEB(WEB),
		.A(A),
		.D(D),
		.BWEB(BWEB),
		.Q(Q)
	);
endmodule
module ram1p1rwbe_64x22 (
	CLK,
	CEB,
	WEB,
	A,
	D,
	BWEB,
	Q
);
	input wire CLK;
	input wire CEB;
	input wire WEB;
	input wire [5:0] A;
	input wire [21:0] D;
	input wire [21:0] BWEB;
	output wire [21:0] Q;
	wire [43:0] Qfull;
	TS1N28HPCPSVTB64X44M4SW sramIP(
		.CLK(CLK),
		.CEB(CEB),
		.WEB(WEB),
		.A(A),
		.D({22'b0000000000000000000000, D[21:0]}),
		.BWEB({22'b0000000000000000000000, BWEB[21:0]}),
		.Q(Qfull)
	);
	assign Q = Qfull[21:0];
endmodule
module ram1p1rwbe_64x44 (
	CLK,
	CEB,
	WEB,
	A,
	D,
	BWEB,
	Q
);
	input wire CLK;
	input wire CEB;
	input wire WEB;
	input wire [5:0] A;
	input wire [43:0] D;
	input wire [43:0] BWEB;
	output wire [43:0] Q;
	TS1N28HPCPSVTB64X44M4SW sramIP(
		.CLK(CLK),
		.CEB(CEB),
		.WEB(WEB),
		.A(A),
		.D(D),
		.BWEB(BWEB),
		.Q(Q)
	);
endmodule
module ram1p1rwe (
	clk,
	ce,
	addr,
	din,
	we,
	dout
);
	parameter USE_SRAM = 0;
	parameter DEPTH = 64;
	parameter WIDTH = 44;
	input wire clk;
	input wire ce;
	input wire [$clog2(DEPTH) - 1:0] addr;
	input wire [WIDTH - 1:0] din;
	input wire we;
	output wire [WIDTH - 1:0] dout;
	generate
		if (((USE_SRAM == 1) & (WIDTH == 128)) & (DEPTH == 64)) begin : genblk1
			localparam [127:0] sv2v_uu_sram1A_ext_BWEB_0 = 1'sb0;
			ram1p1rwbe_64x128 sram1A(
				.CLK(clk),
				.CEB(~ce),
				.WEB(~we),
				.A(addr),
				.D(din),
				.BWEB(sv2v_uu_sram1A_ext_BWEB_0),
				.Q(dout)
			);
		end
		else if (((USE_SRAM == 1) & (WIDTH == 44)) & (DEPTH == 64)) begin : genblk1
			localparam [43:0] sv2v_uu_sram1B_ext_BWEB_0 = 1'sb0;
			ram1p1rwbe_64x44 sram1B(
				.CLK(clk),
				.CEB(~ce),
				.WEB(~we),
				.A(addr),
				.D(din),
				.BWEB(sv2v_uu_sram1B_ext_BWEB_0),
				.Q(dout)
			);
		end
		else if (((USE_SRAM == 1) & (WIDTH == 22)) & (DEPTH == 64)) begin : genblk1
			localparam [21:0] sv2v_uu_sram1_ext_BWEB_0 = 1'sb0;
			ram1p1rwbe_64x22 sram1(
				.CLK(clk),
				.CEB(~ce),
				.WEB(~we),
				.A(addr),
				.D(din),
				.BWEB(sv2v_uu_sram1_ext_BWEB_0),
				.Q(dout)
			);
		end
		else begin : ram
			reg [WIDTH - 1:0] RAM [DEPTH - 1:0];
			wire [$clog2(DEPTH) - 1:0] addrd;
			flopen #(.WIDTH($clog2(DEPTH))) adrreg(
				.clk(clk),
				.en(ce),
				.d(addr),
				.q(addrd)
			);
			assign dout = RAM[addrd];
			always @(posedge clk)
				if (ce & we)
					RAM[addr] <= din;
		end
	endgenerate
endmodule
module ram2p1r1wbe (
	clk,
	ce1,
	ce2,
	ra1,
	wd2,
	wa2,
	we2,
	bwe2,
	rd1
);
	parameter USE_SRAM = 0;
	parameter DEPTH = 1024;
	parameter WIDTH = 68;
	input wire clk;
	input wire ce1;
	input wire ce2;
	input wire [$clog2(DEPTH) - 1:0] ra1;
	input wire [WIDTH - 1:0] wd2;
	input wire [$clog2(DEPTH) - 1:0] wa2;
	input wire we2;
	input wire [(WIDTH - 1) / 8:0] bwe2;
	output wire [WIDTH - 1:0] rd1;
	localparam SRAMWIDTH = 32;
	localparam SRAMNUMSETS = SRAMWIDTH / WIDTH;
	generate
		if (((USE_SRAM == 1) & (WIDTH == 68)) & (DEPTH == 1024)) begin : genblk1
			localparam [67:0] sv2v_uu_memory1_ext_DA_0 = 1'sb0;
			localparam [67:0] sv2v_uu_memory1_ext_BWEBA_0 = 1'sb0;
			localparam [67:0] sv2v_uu_memory1_ext_BWEBB_1 = 1'sb1;
			ram2p1r1wbe_1024x68 memory1(
				.CLKA(clk),
				.CLKB(clk),
				.CEBA(~ce1),
				.CEBB(~ce2),
				.WEBA(1'b0),
				.WEBB(~we2),
				.AA(ra1),
				.AB(wa2),
				.DA(sv2v_uu_memory1_ext_DA_0),
				.DB(wd2),
				.BWEBA(sv2v_uu_memory1_ext_BWEBA_0),
				.BWEBB(sv2v_uu_memory1_ext_BWEBB_1),
				.QA(rd1),
				.QB()
			);
		end
		else if (((USE_SRAM == 1) & (WIDTH == 36)) & (DEPTH == 1024)) begin : genblk1
			localparam [35:0] sv2v_uu_memory1_ext_DA_0 = 1'sb0;
			localparam [35:0] sv2v_uu_memory1_ext_BWEBA_0 = 1'sb0;
			localparam [35:0] sv2v_uu_memory1_ext_BWEBB_1 = 1'sb1;
			ram2p1r1wbe_1024x36 memory1(
				.CLKA(clk),
				.CLKB(clk),
				.CEBA(~ce1),
				.CEBB(~ce2),
				.WEBA(1'b0),
				.WEBB(~we2),
				.AA(ra1),
				.AB(wa2),
				.DA(sv2v_uu_memory1_ext_DA_0),
				.DB(wd2),
				.BWEBA(sv2v_uu_memory1_ext_BWEBA_0),
				.BWEBB(sv2v_uu_memory1_ext_BWEBB_1),
				.QA(rd1),
				.QB()
			);
		end
		else if (((USE_SRAM == 1) & (WIDTH == 2)) & (DEPTH == 1024)) begin : genblk1
			wire [31:0] SRAMReadData;
			wire [31:0] SRAMWriteData;
			wire [31:0] RD1Sets [SRAMNUMSETS - 1:0];
			wire [SRAMNUMSETS - 1:0] SRAMBitMaskPre;
			wire [31:0] SRAMBitMask;
			wire [$clog2(DEPTH) - 1:0] RA1Q;
			onehotdecoder #(.WIDTH($clog2(SRAMNUMSETS))) oh1(
				.bin(wa2[$clog2(SRAMNUMSETS) - 1:0]),
				.decoded(SRAMBitMaskPre)
			);
			genvar _gv_index_11;
			for (_gv_index_11 = 0; _gv_index_11 < SRAMNUMSETS; _gv_index_11 = _gv_index_11 + 1) begin : readdatalinesetsmux
				localparam index = _gv_index_11;
				assign RD1Sets[index] = SRAMReadData[((index * WIDTH) + WIDTH) - 1:index * WIDTH];
				assign SRAMWriteData[(index * 2) + 1:index * 2] = wd2;
				assign SRAMBitMask[(index * 2) + 1:index * 2] = {2 {SRAMBitMaskPre[index]}};
			end
			flopen #(.WIDTH($clog2(DEPTH))) mem_reg1(
				.clk(clk),
				.en(ce1),
				.d(ra1),
				.q(RA1Q)
			);
			assign rd1 = RD1Sets[RA1Q[4:0]];
			localparam [31:0] sv2v_uu_memory2_ext_DA_0 = 1'sb0;
			localparam [31:0] sv2v_uu_memory2_ext_BWEBA_0 = 1'sb0;
			ram2p1r1wbe_64x32 memory2(
				.CLKA(clk),
				.CLKB(clk),
				.CEBA(~ce1),
				.CEBB(~ce2),
				.WEBA(1'b0),
				.WEBB(~we2),
				.AA(ra1[$clog2(DEPTH) - 1:$clog2(SRAMNUMSETS)]),
				.AB(wa2[$clog2(DEPTH) - 1:$clog2(SRAMNUMSETS)]),
				.DA(sv2v_uu_memory2_ext_DA_0),
				.DB(SRAMWriteData),
				.BWEBA(sv2v_uu_memory2_ext_BWEBA_0),
				.BWEBB(SRAMBitMask),
				.QA(SRAMReadData),
				.QB()
			);
		end
		else begin : ram
			reg [WIDTH - 1:0] RAM [DEPTH - 1:0];
			wire [$clog2(DEPTH) - 1:0] ra1d;
			flopen #(.WIDTH($clog2(DEPTH))) adrreg(
				.clk(clk),
				.en(ce1),
				.d(ra1),
				.q(ra1d)
			);
			assign rd1 = RAM[ra1d];
			if (WIDTH >= 8) begin : genblk1
				integer i;
				always @(posedge clk)
					if (ce2 & we2) begin
						for (i = 0; i < (WIDTH / 8); i = i + 1)
							if (bwe2[i])
								RAM[wa2][i * 8+:8] <= wd2[i * 8+:8];
					end
			end
			if ((WIDTH % 8) != 0) begin : genblk2
				always @(posedge clk)
					if ((ce2 & we2) & bwe2[WIDTH / 8])
						RAM[wa2][WIDTH - 1:WIDTH - (WIDTH % 8)] <= wd2[WIDTH - 1:WIDTH - (WIDTH % 8)];
			end
		end
	endgenerate
endmodule
module ram2p1r1wbe_1024x36 (
	CLKA,
	CLKB,
	CEBA,
	CEBB,
	WEBA,
	WEBB,
	AA,
	AB,
	DA,
	DB,
	BWEBA,
	BWEBB,
	QA,
	QB
);
	input wire CLKA;
	input wire CLKB;
	input wire CEBA;
	input wire CEBB;
	input wire WEBA;
	input wire WEBB;
	input wire [9:0] AA;
	input wire [9:0] AB;
	input wire [35:0] DA;
	input wire [35:0] DB;
	input wire [35:0] BWEBA;
	input wire [35:0] BWEBB;
	output wire [35:0] QA;
	output wire [35:0] QB;
	wire [67:0] QAfull;
	wire [67:0] QBfull;
	TSDN28HPCPA1024X68M4MW sramIP(
		.CLKA(CLKA),
		.CLKB(CLKB),
		.CEBA(CEBA),
		.CEBB(CEBB),
		.WEBA(WEBA),
		.WEBB(WEBB),
		.AA(AA),
		.AB(AB),
		.DA({32'b00000000000000000000000000000000, DA[35:0]}),
		.DB({32'b00000000000000000000000000000000, DB[35:0]}),
		.BWEBA({32'b00000000000000000000000000000000, BWEBA[35:0]}),
		.BWEBB({32'b00000000000000000000000000000000, BWEBB[35:0]}),
		.QA(QAfull),
		.QB(QBfull)
	);
	assign QA = QAfull[35:0];
	assign QB = QBfull[35:0];
endmodule
module ram2p1r1wbe_1024x68 (
	CLKA,
	CLKB,
	CEBA,
	CEBB,
	WEBA,
	WEBB,
	AA,
	AB,
	DA,
	DB,
	BWEBA,
	BWEBB,
	QA,
	QB
);
	input wire CLKA;
	input wire CLKB;
	input wire CEBA;
	input wire CEBB;
	input wire WEBA;
	input wire WEBB;
	input wire [9:0] AA;
	input wire [9:0] AB;
	input wire [67:0] DA;
	input wire [67:0] DB;
	input wire [67:0] BWEBA;
	input wire [67:0] BWEBB;
	output wire [67:0] QA;
	output wire [67:0] QB;
	TSDN28HPCPA1024X68M4MW sramIP(
		.CLKA(CLKA),
		.CLKB(CLKB),
		.CEBA(CEBA),
		.CEBB(CEBB),
		.WEBA(WEBA),
		.WEBB(WEBB),
		.AA(AA),
		.AB(AB),
		.DA(DA),
		.DB(DB),
		.BWEBA(BWEBA),
		.BWEBB(BWEBB),
		.QA(QA),
		.QB(QB)
	);
endmodule
module ram2p1r1wbe_128x64 (
	CLKA,
	CLKB,
	CEBA,
	CEBB,
	WEBA,
	WEBB,
	AA,
	AB,
	DA,
	DB,
	BWEBA,
	BWEBB,
	QA,
	QB
);
	input wire CLKA;
	input wire CLKB;
	input wire CEBA;
	input wire CEBB;
	input wire WEBA;
	input wire WEBB;
	input wire [6:0] AA;
	input wire [6:0] AB;
	input wire [63:0] DA;
	input wire [63:0] DB;
	input wire [63:0] BWEBA;
	input wire [63:0] BWEBB;
	output wire [63:0] QA;
	output wire [63:0] QB;
	TSDN28HPCPA128X64M4FW sramIP(
		.CLKA(CLKA),
		.CLKB(CLKB),
		.CEBA(CEBA),
		.CEBB(CEBB),
		.WEBA(WEBA),
		.WEBB(WEBB),
		.AA(AA),
		.AB(AB),
		.DA(DA),
		.DB(DB),
		.BWEBA(BWEBA),
		.BWEBB(BWEBB),
		.QA(QA),
		.QB(QB)
	);
endmodule
module ram2p1r1wbe_2048x64 (
	CLKA,
	CLKB,
	CEBA,
	CEBB,
	WEBA,
	WEBB,
	AA,
	AB,
	DA,
	DB,
	BWEBA,
	BWEBB,
	QA,
	QB
);
	input wire CLKA;
	input wire CLKB;
	input wire CEBA;
	input wire CEBB;
	input wire WEBA;
	input wire WEBB;
	input wire [8:0] AA;
	input wire [8:0] AB;
	input wire [63:0] DA;
	input wire [63:0] DB;
	input wire [63:0] BWEBA;
	input wire [63:0] BWEBB;
	output wire [63:0] QA;
	output wire [63:0] QB;
	TSDN28HPCPA2048X64MMFW sramIP(
		.CLKA(CLKA),
		.CLKB(CLKB),
		.CEBA(CEBA),
		.CEBB(CEBB),
		.WEBA(WEBA),
		.WEBB(WEBB),
		.AA(AA),
		.AB(AB),
		.DA(DA),
		.DB(DB),
		.BWEBA(BWEBA),
		.BWEBB(BWEBB),
		.QA(QA),
		.QB(QB)
	);
endmodule
module ram2p1r1wbe_64x32 (
	CLKA,
	CLKB,
	CEBA,
	CEBB,
	WEBA,
	WEBB,
	AA,
	AB,
	DA,
	DB,
	BWEBA,
	BWEBB,
	QA,
	QB
);
	input wire CLKA;
	input wire CLKB;
	input wire CEBA;
	input wire CEBB;
	input wire WEBA;
	input wire WEBB;
	input wire [5:0] AA;
	input wire [5:0] AB;
	input wire [31:0] DA;
	input wire [31:0] DB;
	input wire [31:0] BWEBA;
	input wire [31:0] BWEBB;
	output wire [31:0] QA;
	output wire [31:0] QB;
	TSDN28HPCPA64X32M4MW sramIP(
		.CLKA(CLKA),
		.CLKB(CLKB),
		.CEBA(CEBA),
		.CEBB(CEBB),
		.WEBA(WEBA),
		.WEBB(WEBB),
		.AA(AA),
		.AB(AB),
		.DA(DA),
		.DB(DB),
		.BWEBA(BWEBA),
		.BWEBB(BWEBB),
		.QA(QA),
		.QB(QB)
	);
endmodule
module rom1p1r (
	clk,
	ce,
	addr,
	dout
);
	parameter ADDR_WIDTH = 8;
	parameter DATA_WIDTH = 32;
	parameter PRELOAD_ENABLED = 0;
	input wire clk;
	input wire ce;
	input wire [ADDR_WIDTH - 1:0] addr;
	output reg [DATA_WIDTH - 1:0] dout;
	reg [DATA_WIDTH - 1:0] ROM [(2 ** ADDR_WIDTH) - 1:0];
	initial if (PRELOAD_ENABLED) begin
		if (DATA_WIDTH == 64)
			$readmemh({"$WALLY/fpga/src/boot.mem"}, ROM, 0);
		else
			ROM[0] = 'h2197;
	end
	always @(posedge clk)
		if (ce)
			dout <= ROM[addr];
endmodule
module rom1p1r_128x32 (
	CLK,
	CEB,
	A,
	Q
);
	input wire CLK;
	input wire CEB;
	input wire [6:0] A;
	output wire [31:0] Q;
	generic64x128ROM sramIP(
		.CLK(CLK),
		.CEB(CEB),
		.A(A),
		.Q(Q)
	);
endmodule
module rom1p1r_128x64 (
	CLK,
	CEB,
	A,
	Q
);
	input wire CLK;
	input wire CEB;
	input wire [6:0] A;
	output wire [63:0] Q;
	ts3n28hpcpa128x64m8m romIP(
		.CLK(CLK),
		.CEB(CEB),
		.A(A),
		.Q(Q)
	);
endmodule
module aes32d (
	SboxIn,
	finalround,
	result
);
	input wire [7:0] SboxIn;
	input wire finalround;
	output wire [31:0] result;
	wire [7:0] SboxOut;
	wire [31:0] so;
	wire [31:0] mixed;
	aesinvsbox8 inv_sbox(
		.a(SboxIn),
		.y(SboxOut)
	);
	aesinvmixcolumns8 mix(
		.a(SboxOut),
		.y(mixed)
	);
	assign so = {24'h000000, SboxOut};
	mux2 #(.WIDTH(32)) rmux(
		.d0(mixed),
		.d1(so),
		.s(finalround),
		.y(result)
	);
endmodule
module aes32e (
	SboxIn,
	finalround,
	result
);
	input wire [7:0] SboxIn;
	input wire finalround;
	output wire [31:0] result;
	wire [7:0] SboxOut;
	wire [31:0] so;
	wire [31:0] mixed;
	aessbox8 sbox(
		.a(SboxIn),
		.y(SboxOut)
	);
	assign so = {24'h000000, SboxOut};
	aesmixcolumns32 mb(
		.a(so),
		.y(mixed)
	);
	mux2 #(.WIDTH(32)) rmux(
		.d0(mixed),
		.d1(so),
		.s(finalround),
		.y(result)
	);
endmodule
module aes64d (
	rs1,
	rs2,
	finalround,
	aes64im,
	result
);
	input wire [63:0] rs1;
	input wire [63:0] rs2;
	input wire finalround;
	input wire aes64im;
	output wire [63:0] result;
	wire [63:0] ShiftRowsOut;
	wire [63:0] SboxOut;
	wire [63:0] MixcolsIn;
	wire [63:0] MixcolsOut;
	aesinvshiftrows64 srow(
		.a({rs2, rs1}),
		.y(ShiftRowsOut)
	);
	aesinvsbox64 invsbox(
		.a(ShiftRowsOut),
		.y(SboxOut)
	);
	mux2 #(.WIDTH(64)) mixcolmux(
		.d0(SboxOut),
		.d1(rs1),
		.s(aes64im),
		.y(MixcolsIn)
	);
	aesinvmixcolumns32 invmw0(
		.a(MixcolsIn[31:0]),
		.y(MixcolsOut[31:0])
	);
	aesinvmixcolumns32 invmw1(
		.a(MixcolsIn[63:32]),
		.y(MixcolsOut[63:32])
	);
	mux2 #(.WIDTH(64)) resultmux(
		.d0(MixcolsOut),
		.d1(SboxOut),
		.s(finalround),
		.y(result)
	);
endmodule
module aes64e (
	rs1,
	rs2,
	finalround,
	Sbox0Out,
	SboxEIn,
	result
);
	input wire [63:0] rs1;
	input wire [63:0] rs2;
	input wire finalround;
	input wire [31:0] Sbox0Out;
	output wire [31:0] SboxEIn;
	output wire [63:0] result;
	wire [63:0] ShiftRowsOut;
	wire [63:0] SboxOut;
	wire [63:0] MixcolsOut;
	aesshiftrows64 srow(
		.a({rs2, rs1}),
		.y(ShiftRowsOut)
	);
	assign SboxEIn = ShiftRowsOut[31:0];
	assign SboxOut[31:0] = Sbox0Out;
	aessbox32 sbox1(
		.a(ShiftRowsOut[63:32]),
		.y(SboxOut[63:32])
	);
	aesmixcolumns32 mw0(
		.a(SboxOut[31:0]),
		.y(MixcolsOut[31:0])
	);
	aesmixcolumns32 mw1(
		.a(SboxOut[63:32]),
		.y(MixcolsOut[63:32])
	);
	mux2 #(.WIDTH(64)) resultmux(
		.d0(MixcolsOut),
		.d1(SboxOut),
		.s(finalround),
		.y(result)
	);
endmodule
module aes64ks1i (
	round,
	rs1,
	Sbox0Out,
	SboxKIn,
	result
);
	input wire [3:0] round;
	input wire [63:32] rs1;
	input wire [31:0] Sbox0Out;
	output wire [31:0] SboxKIn;
	output wire [63:0] result;
	wire finalround;
	wire [31:0] rcon;
	wire [31:0] rs1Rotate;
	rconlut32 rc(
		.rd(round),
		.rcon(rcon)
	);
	assign rs1Rotate = {rs1[39:32], rs1[63:40]};
	assign finalround = round == 4'b1010;
	assign SboxKIn = (finalround ? rs1[63:32] : rs1Rotate);
	assign result[31:0] = Sbox0Out ^ rcon;
	assign result[63:32] = Sbox0Out ^ rcon;
endmodule
module aes64ks2 (
	rs2,
	rs1,
	result
);
	input wire [63:0] rs2;
	input wire [63:32] rs1;
	output wire [63:0] result;
	wire [31:0] w0;
	wire [31:0] w1;
	assign w0 = rs1[63:32] ^ rs2[31:0];
	assign w1 = w0 ^ rs2[63:32];
	assign result = {w1, w0};
endmodule
module aesinvmixcolumns32 (
	a,
	y
);
	input wire [31:0] a;
	output wire [31:0] y;
	wire [7:0] a0;
	wire [7:0] a1;
	wire [7:0] a2;
	wire [7:0] a3;
	wire [7:0] temp;
	wire [10:0] xor0;
	wire [10:0] xor1;
	wire [10:0] xor2;
	wire [10:0] xor3;
	assign {a0, a1, a2, a3} = a;
	assign temp = ((a0 ^ a1) ^ a2) ^ a3;
	assign xor0 = ((({temp, 3'b000} ^ {1'b0, a3 ^ a1, 2'b00}) ^ {2'b00, a3 ^ a2, 1'b0}) ^ {3'b000, temp}) ^ {3'b000, a3};
	assign xor1 = ((({temp, 3'b000} ^ {1'b0, a2 ^ a0, 2'b00}) ^ {2'b00, a2 ^ a1, 1'b0}) ^ {3'b000, temp}) ^ {3'b000, a2};
	assign xor2 = ((({temp, 3'b000} ^ {1'b0, a1 ^ a3, 2'b00}) ^ {2'b00, a1 ^ a0, 1'b0}) ^ {3'b000, temp}) ^ {3'b000, a1};
	assign xor3 = ((({temp, 3'b000} ^ {1'b0, a0 ^ a2, 2'b00}) ^ {2'b00, a0 ^ a3, 1'b0}) ^ {3'b000, temp}) ^ {3'b000, a0};
	galoismultinverse8 gm0(
		.a(xor0),
		.y(y[7:0])
	);
	galoismultinverse8 gm1(
		.a(xor1),
		.y(y[15:8])
	);
	galoismultinverse8 gm2(
		.a(xor2),
		.y(y[23:16])
	);
	galoismultinverse8 gm3(
		.a(xor3),
		.y(y[31:24])
	);
endmodule
module aesinvmixcolumns8 (
	a,
	y
);
	input wire [7:0] a;
	output wire [31:0] y;
	wire [10:0] t;
	wire [10:0] x0;
	wire [10:0] x1;
	wire [10:0] x2;
	wire [10:0] x3;
	assign t = {a, 3'b000} ^ {3'b000, a};
	assign x0 = ({a, 3'b000} ^ {1'b0, a, 2'b00}) ^ {2'b00, a, 1'b0};
	assign x1 = t;
	assign x2 = t ^ {1'b0, a, 2'b00};
	assign x3 = t ^ {2'b00, a, 1'b0};
	galoismultinverse8 gm0(
		.a(x0),
		.y(y[7:0])
	);
	galoismultinverse8 gm1(
		.a(x1),
		.y(y[15:8])
	);
	galoismultinverse8 gm2(
		.a(x2),
		.y(y[23:16])
	);
	galoismultinverse8 gm3(
		.a(x3),
		.y(y[31:24])
	);
endmodule
module aesinvsbox64 (
	a,
	y
);
	input wire [63:0] a;
	output wire [63:0] y;
	aesinvsbox8 sbox0(
		.a(a[7:0]),
		.y(y[7:0])
	);
	aesinvsbox8 sbox1(
		.a(a[15:8]),
		.y(y[15:8])
	);
	aesinvsbox8 sbox2(
		.a(a[23:16]),
		.y(y[23:16])
	);
	aesinvsbox8 sbox3(
		.a(a[31:24]),
		.y(y[31:24])
	);
	aesinvsbox8 sbox4(
		.a(a[39:32]),
		.y(y[39:32])
	);
	aesinvsbox8 sbox5(
		.a(a[47:40]),
		.y(y[47:40])
	);
	aesinvsbox8 sbox6(
		.a(a[55:48]),
		.y(y[55:48])
	);
	aesinvsbox8 sbox7(
		.a(a[63:56]),
		.y(y[63:56])
	);
endmodule
module aesinvsbox8 (
	a,
	y
);
	reg _sv2v_0;
	input wire [7:0] a;
	output reg [7:0] y;
	always @(*) begin
		if (_sv2v_0)
			;
		case (a)
			8'h00: y = 8'h52;
			8'h01: y = 8'h09;
			8'h02: y = 8'h6a;
			8'h03: y = 8'hd5;
			8'h04: y = 8'h30;
			8'h05: y = 8'h36;
			8'h06: y = 8'ha5;
			8'h07: y = 8'h38;
			8'h08: y = 8'hbf;
			8'h09: y = 8'h40;
			8'h0a: y = 8'ha3;
			8'h0b: y = 8'h9e;
			8'h0c: y = 8'h81;
			8'h0d: y = 8'hf3;
			8'h0e: y = 8'hd7;
			8'h0f: y = 8'hfb;
			8'h10: y = 8'h7c;
			8'h11: y = 8'he3;
			8'h12: y = 8'h39;
			8'h13: y = 8'h82;
			8'h14: y = 8'h9b;
			8'h15: y = 8'h2f;
			8'h16: y = 8'hff;
			8'h17: y = 8'h87;
			8'h18: y = 8'h34;
			8'h19: y = 8'h8e;
			8'h1a: y = 8'h43;
			8'h1b: y = 8'h44;
			8'h1c: y = 8'hc4;
			8'h1d: y = 8'hde;
			8'h1e: y = 8'he9;
			8'h1f: y = 8'hcb;
			8'h20: y = 8'h54;
			8'h21: y = 8'h7b;
			8'h22: y = 8'h94;
			8'h23: y = 8'h32;
			8'h24: y = 8'ha6;
			8'h25: y = 8'hc2;
			8'h26: y = 8'h23;
			8'h27: y = 8'h3d;
			8'h28: y = 8'hee;
			8'h29: y = 8'h4c;
			8'h2a: y = 8'h95;
			8'h2b: y = 8'h0b;
			8'h2c: y = 8'h42;
			8'h2d: y = 8'hfa;
			8'h2e: y = 8'hc3;
			8'h2f: y = 8'h4e;
			8'h30: y = 8'h08;
			8'h31: y = 8'h2e;
			8'h32: y = 8'ha1;
			8'h33: y = 8'h66;
			8'h34: y = 8'h28;
			8'h35: y = 8'hd9;
			8'h36: y = 8'h24;
			8'h37: y = 8'hb2;
			8'h38: y = 8'h76;
			8'h39: y = 8'h5b;
			8'h3a: y = 8'ha2;
			8'h3b: y = 8'h49;
			8'h3c: y = 8'h6d;
			8'h3d: y = 8'h8b;
			8'h3e: y = 8'hd1;
			8'h3f: y = 8'h25;
			8'h40: y = 8'h72;
			8'h41: y = 8'hf8;
			8'h42: y = 8'hf6;
			8'h43: y = 8'h64;
			8'h44: y = 8'h86;
			8'h45: y = 8'h68;
			8'h46: y = 8'h98;
			8'h47: y = 8'h16;
			8'h48: y = 8'hd4;
			8'h49: y = 8'ha4;
			8'h4a: y = 8'h5c;
			8'h4b: y = 8'hcc;
			8'h4c: y = 8'h5d;
			8'h4d: y = 8'h65;
			8'h4e: y = 8'hb6;
			8'h4f: y = 8'h92;
			8'h50: y = 8'h6c;
			8'h51: y = 8'h70;
			8'h52: y = 8'h48;
			8'h53: y = 8'h50;
			8'h54: y = 8'hfd;
			8'h55: y = 8'hed;
			8'h56: y = 8'hb9;
			8'h57: y = 8'hda;
			8'h58: y = 8'h5e;
			8'h59: y = 8'h15;
			8'h5a: y = 8'h46;
			8'h5b: y = 8'h57;
			8'h5c: y = 8'ha7;
			8'h5d: y = 8'h8d;
			8'h5e: y = 8'h9d;
			8'h5f: y = 8'h84;
			8'h60: y = 8'h90;
			8'h61: y = 8'hd8;
			8'h62: y = 8'hab;
			8'h63: y = 8'h00;
			8'h64: y = 8'h8c;
			8'h65: y = 8'hbc;
			8'h66: y = 8'hd3;
			8'h67: y = 8'h0a;
			8'h68: y = 8'hf7;
			8'h69: y = 8'he4;
			8'h6a: y = 8'h58;
			8'h6b: y = 8'h05;
			8'h6c: y = 8'hb8;
			8'h6d: y = 8'hb3;
			8'h6e: y = 8'h45;
			8'h6f: y = 8'h06;
			8'h70: y = 8'hd0;
			8'h71: y = 8'h2c;
			8'h72: y = 8'h1e;
			8'h73: y = 8'h8f;
			8'h74: y = 8'hca;
			8'h75: y = 8'h3f;
			8'h76: y = 8'h0f;
			8'h77: y = 8'h02;
			8'h78: y = 8'hc1;
			8'h79: y = 8'haf;
			8'h7a: y = 8'hbd;
			8'h7b: y = 8'h03;
			8'h7c: y = 8'h01;
			8'h7d: y = 8'h13;
			8'h7e: y = 8'h8a;
			8'h7f: y = 8'h6b;
			8'h80: y = 8'h3a;
			8'h81: y = 8'h91;
			8'h82: y = 8'h11;
			8'h83: y = 8'h41;
			8'h84: y = 8'h4f;
			8'h85: y = 8'h67;
			8'h86: y = 8'hdc;
			8'h87: y = 8'hea;
			8'h88: y = 8'h97;
			8'h89: y = 8'hf2;
			8'h8a: y = 8'hcf;
			8'h8b: y = 8'hce;
			8'h8c: y = 8'hf0;
			8'h8d: y = 8'hb4;
			8'h8e: y = 8'he6;
			8'h8f: y = 8'h73;
			8'h90: y = 8'h96;
			8'h91: y = 8'hac;
			8'h92: y = 8'h74;
			8'h93: y = 8'h22;
			8'h94: y = 8'he7;
			8'h95: y = 8'had;
			8'h96: y = 8'h35;
			8'h97: y = 8'h85;
			8'h98: y = 8'he2;
			8'h99: y = 8'hf9;
			8'h9a: y = 8'h37;
			8'h9b: y = 8'he8;
			8'h9c: y = 8'h1c;
			8'h9d: y = 8'h75;
			8'h9e: y = 8'hdf;
			8'h9f: y = 8'h6e;
			8'ha0: y = 8'h47;
			8'ha1: y = 8'hf1;
			8'ha2: y = 8'h1a;
			8'ha3: y = 8'h71;
			8'ha4: y = 8'h1d;
			8'ha5: y = 8'h29;
			8'ha6: y = 8'hc5;
			8'ha7: y = 8'h89;
			8'ha8: y = 8'h6f;
			8'ha9: y = 8'hb7;
			8'haa: y = 8'h62;
			8'hab: y = 8'h0e;
			8'hac: y = 8'haa;
			8'had: y = 8'h18;
			8'hae: y = 8'hbe;
			8'haf: y = 8'h1b;
			8'hb0: y = 8'hfc;
			8'hb1: y = 8'h56;
			8'hb2: y = 8'h3e;
			8'hb3: y = 8'h4b;
			8'hb4: y = 8'hc6;
			8'hb5: y = 8'hd2;
			8'hb6: y = 8'h79;
			8'hb7: y = 8'h20;
			8'hb8: y = 8'h9a;
			8'hb9: y = 8'hdb;
			8'hba: y = 8'hc0;
			8'hbb: y = 8'hfe;
			8'hbc: y = 8'h78;
			8'hbd: y = 8'hcd;
			8'hbe: y = 8'h5a;
			8'hbf: y = 8'hf4;
			8'hc0: y = 8'h1f;
			8'hc1: y = 8'hdd;
			8'hc2: y = 8'ha8;
			8'hc3: y = 8'h33;
			8'hc4: y = 8'h88;
			8'hc5: y = 8'h07;
			8'hc6: y = 8'hc7;
			8'hc7: y = 8'h31;
			8'hc8: y = 8'hb1;
			8'hc9: y = 8'h12;
			8'hca: y = 8'h10;
			8'hcb: y = 8'h59;
			8'hcc: y = 8'h27;
			8'hcd: y = 8'h80;
			8'hce: y = 8'hec;
			8'hcf: y = 8'h5f;
			8'hd0: y = 8'h60;
			8'hd1: y = 8'h51;
			8'hd2: y = 8'h7f;
			8'hd3: y = 8'ha9;
			8'hd4: y = 8'h19;
			8'hd5: y = 8'hb5;
			8'hd6: y = 8'h4a;
			8'hd7: y = 8'h0d;
			8'hd8: y = 8'h2d;
			8'hd9: y = 8'he5;
			8'hda: y = 8'h7a;
			8'hdb: y = 8'h9f;
			8'hdc: y = 8'h93;
			8'hdd: y = 8'hc9;
			8'hde: y = 8'h9c;
			8'hdf: y = 8'hef;
			8'he0: y = 8'ha0;
			8'he1: y = 8'he0;
			8'he2: y = 8'h3b;
			8'he3: y = 8'h4d;
			8'he4: y = 8'hae;
			8'he5: y = 8'h2a;
			8'he6: y = 8'hf5;
			8'he7: y = 8'hb0;
			8'he8: y = 8'hc8;
			8'he9: y = 8'heb;
			8'hea: y = 8'hbb;
			8'heb: y = 8'h3c;
			8'hec: y = 8'h83;
			8'hed: y = 8'h53;
			8'hee: y = 8'h99;
			8'hef: y = 8'h61;
			8'hf0: y = 8'h17;
			8'hf1: y = 8'h2b;
			8'hf2: y = 8'h04;
			8'hf3: y = 8'h7e;
			8'hf4: y = 8'hba;
			8'hf5: y = 8'h77;
			8'hf6: y = 8'hd6;
			8'hf7: y = 8'h26;
			8'hf8: y = 8'he1;
			8'hf9: y = 8'h69;
			8'hfa: y = 8'h14;
			8'hfb: y = 8'h63;
			8'hfc: y = 8'h55;
			8'hfd: y = 8'h21;
			8'hfe: y = 8'h0c;
			8'hff: y = 8'h7d;
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
module aesinvshiftrows64 (
	a,
	y
);
	input wire [127:0] a;
	output wire [63:0] y;
	assign y = {a[95:88], a[119:112], a[15:8], a[39:32], a[63:56], a[87:80], a[111:104], a[7:0]};
endmodule
module aesmixcolumns32 (
	a,
	y
);
	input wire [31:0] a;
	output wire [31:0] y;
	wire [7:0] a0;
	wire [7:0] a1;
	wire [7:0] a2;
	wire [7:0] a3;
	wire [7:0] y0;
	wire [7:0] y1;
	wire [7:0] y2;
	wire [7:0] y3;
	wire [7:0] t0;
	wire [7:0] t1;
	wire [7:0] t2;
	wire [7:0] t3;
	wire [7:0] temp;
	assign {a0, a1, a2, a3} = a;
	assign temp = ((a0 ^ a1) ^ a2) ^ a3;
	galoismultforward8 gm0(
		.a(a0 ^ a1),
		.y(t0)
	);
	galoismultforward8 gm1(
		.a(a1 ^ a2),
		.y(t1)
	);
	galoismultforward8 gm2(
		.a(a2 ^ a3),
		.y(t2)
	);
	galoismultforward8 gm3(
		.a(a3 ^ a0),
		.y(t3)
	);
	assign y0 = (a0 ^ temp) ^ t3;
	assign y1 = (a1 ^ temp) ^ t0;
	assign y2 = (a2 ^ temp) ^ t1;
	assign y3 = (a3 ^ temp) ^ t2;
	assign y = {y0, y1, y2, y3};
endmodule
module aesmixcolumns8 (
	a,
	y
);
	input wire [7:0] a;
	output wire [31:0] y;
	wire [7:0] xa;
	wire [7:0] xapa;
	galoismultforward8 gm(
		.a(a),
		.y(xa)
	);
	assign xapa = a ^ xa;
	assign y = {xapa, a, a, xa};
endmodule
module aessbox32 (
	a,
	y
);
	input wire [31:0] a;
	output wire [31:0] y;
	aessbox8 sbox0(
		.a(a[7:0]),
		.y(y[7:0])
	);
	aessbox8 sbox1(
		.a(a[15:8]),
		.y(y[15:8])
	);
	aessbox8 sbox2(
		.a(a[23:16]),
		.y(y[23:16])
	);
	aessbox8 sbox3(
		.a(a[31:24]),
		.y(y[31:24])
	);
endmodule
module aessbox8 (
	a,
	y
);
	reg _sv2v_0;
	input wire [7:0] a;
	output reg [7:0] y;
	always @(*) begin
		if (_sv2v_0)
			;
		case (a)
			8'h00: y = 8'h63;
			8'h01: y = 8'h7c;
			8'h02: y = 8'h77;
			8'h03: y = 8'h7b;
			8'h04: y = 8'hf2;
			8'h05: y = 8'h6b;
			8'h06: y = 8'h6f;
			8'h07: y = 8'hc5;
			8'h08: y = 8'h30;
			8'h09: y = 8'h01;
			8'h0a: y = 8'h67;
			8'h0b: y = 8'h2b;
			8'h0c: y = 8'hfe;
			8'h0d: y = 8'hd7;
			8'h0e: y = 8'hab;
			8'h0f: y = 8'h76;
			8'h10: y = 8'hca;
			8'h11: y = 8'h82;
			8'h12: y = 8'hc9;
			8'h13: y = 8'h7d;
			8'h14: y = 8'hfa;
			8'h15: y = 8'h59;
			8'h16: y = 8'h47;
			8'h17: y = 8'hf0;
			8'h18: y = 8'had;
			8'h19: y = 8'hd4;
			8'h1a: y = 8'ha2;
			8'h1b: y = 8'haf;
			8'h1c: y = 8'h9c;
			8'h1d: y = 8'ha4;
			8'h1e: y = 8'h72;
			8'h1f: y = 8'hc0;
			8'h20: y = 8'hb7;
			8'h21: y = 8'hfd;
			8'h22: y = 8'h93;
			8'h23: y = 8'h26;
			8'h24: y = 8'h36;
			8'h25: y = 8'h3f;
			8'h26: y = 8'hf7;
			8'h27: y = 8'hcc;
			8'h28: y = 8'h34;
			8'h29: y = 8'ha5;
			8'h2a: y = 8'he5;
			8'h2b: y = 8'hf1;
			8'h2c: y = 8'h71;
			8'h2d: y = 8'hd8;
			8'h2e: y = 8'h31;
			8'h2f: y = 8'h15;
			8'h30: y = 8'h04;
			8'h31: y = 8'hc7;
			8'h32: y = 8'h23;
			8'h33: y = 8'hc3;
			8'h34: y = 8'h18;
			8'h35: y = 8'h96;
			8'h36: y = 8'h05;
			8'h37: y = 8'h9a;
			8'h38: y = 8'h07;
			8'h39: y = 8'h12;
			8'h3a: y = 8'h80;
			8'h3b: y = 8'he2;
			8'h3c: y = 8'heb;
			8'h3d: y = 8'h27;
			8'h3e: y = 8'hb2;
			8'h3f: y = 8'h75;
			8'h40: y = 8'h09;
			8'h41: y = 8'h83;
			8'h42: y = 8'h2c;
			8'h43: y = 8'h1a;
			8'h44: y = 8'h1b;
			8'h45: y = 8'h6e;
			8'h46: y = 8'h5a;
			8'h47: y = 8'ha0;
			8'h48: y = 8'h52;
			8'h49: y = 8'h3b;
			8'h4a: y = 8'hd6;
			8'h4b: y = 8'hb3;
			8'h4c: y = 8'h29;
			8'h4d: y = 8'he3;
			8'h4e: y = 8'h2f;
			8'h4f: y = 8'h84;
			8'h50: y = 8'h53;
			8'h51: y = 8'hd1;
			8'h52: y = 8'h00;
			8'h53: y = 8'hed;
			8'h54: y = 8'h20;
			8'h55: y = 8'hfc;
			8'h56: y = 8'hb1;
			8'h57: y = 8'h5b;
			8'h58: y = 8'h6a;
			8'h59: y = 8'hcb;
			8'h5a: y = 8'hbe;
			8'h5b: y = 8'h39;
			8'h5c: y = 8'h4a;
			8'h5d: y = 8'h4c;
			8'h5e: y = 8'h58;
			8'h5f: y = 8'hcf;
			8'h60: y = 8'hd0;
			8'h61: y = 8'hef;
			8'h62: y = 8'haa;
			8'h63: y = 8'hfb;
			8'h64: y = 8'h43;
			8'h65: y = 8'h4d;
			8'h66: y = 8'h33;
			8'h67: y = 8'h85;
			8'h68: y = 8'h45;
			8'h69: y = 8'hf9;
			8'h6a: y = 8'h02;
			8'h6b: y = 8'h7f;
			8'h6c: y = 8'h50;
			8'h6d: y = 8'h3c;
			8'h6e: y = 8'h9f;
			8'h6f: y = 8'ha8;
			8'h70: y = 8'h51;
			8'h71: y = 8'ha3;
			8'h72: y = 8'h40;
			8'h73: y = 8'h8f;
			8'h74: y = 8'h92;
			8'h75: y = 8'h9d;
			8'h76: y = 8'h38;
			8'h77: y = 8'hf5;
			8'h78: y = 8'hbc;
			8'h79: y = 8'hb6;
			8'h7a: y = 8'hda;
			8'h7b: y = 8'h21;
			8'h7c: y = 8'h10;
			8'h7d: y = 8'hff;
			8'h7e: y = 8'hf3;
			8'h7f: y = 8'hd2;
			8'h80: y = 8'hcd;
			8'h81: y = 8'h0c;
			8'h82: y = 8'h13;
			8'h83: y = 8'hec;
			8'h84: y = 8'h5f;
			8'h85: y = 8'h97;
			8'h86: y = 8'h44;
			8'h87: y = 8'h17;
			8'h88: y = 8'hc4;
			8'h89: y = 8'ha7;
			8'h8a: y = 8'h7e;
			8'h8b: y = 8'h3d;
			8'h8c: y = 8'h64;
			8'h8d: y = 8'h5d;
			8'h8e: y = 8'h19;
			8'h8f: y = 8'h73;
			8'h90: y = 8'h60;
			8'h91: y = 8'h81;
			8'h92: y = 8'h4f;
			8'h93: y = 8'hdc;
			8'h94: y = 8'h22;
			8'h95: y = 8'h2a;
			8'h96: y = 8'h90;
			8'h97: y = 8'h88;
			8'h98: y = 8'h46;
			8'h99: y = 8'hee;
			8'h9a: y = 8'hb8;
			8'h9b: y = 8'h14;
			8'h9c: y = 8'hde;
			8'h9d: y = 8'h5e;
			8'h9e: y = 8'h0b;
			8'h9f: y = 8'hdb;
			8'ha0: y = 8'he0;
			8'ha1: y = 8'h32;
			8'ha2: y = 8'h3a;
			8'ha3: y = 8'h0a;
			8'ha4: y = 8'h49;
			8'ha5: y = 8'h06;
			8'ha6: y = 8'h24;
			8'ha7: y = 8'h5c;
			8'ha8: y = 8'hc2;
			8'ha9: y = 8'hd3;
			8'haa: y = 8'hac;
			8'hab: y = 8'h62;
			8'hac: y = 8'h91;
			8'had: y = 8'h95;
			8'hae: y = 8'he4;
			8'haf: y = 8'h79;
			8'hb0: y = 8'he7;
			8'hb1: y = 8'hc8;
			8'hb2: y = 8'h37;
			8'hb3: y = 8'h6d;
			8'hb4: y = 8'h8d;
			8'hb5: y = 8'hd5;
			8'hb6: y = 8'h4e;
			8'hb7: y = 8'ha9;
			8'hb8: y = 8'h6c;
			8'hb9: y = 8'h56;
			8'hba: y = 8'hf4;
			8'hbb: y = 8'hea;
			8'hbc: y = 8'h65;
			8'hbd: y = 8'h7a;
			8'hbe: y = 8'hae;
			8'hbf: y = 8'h08;
			8'hc0: y = 8'hba;
			8'hc1: y = 8'h78;
			8'hc2: y = 8'h25;
			8'hc3: y = 8'h2e;
			8'hc4: y = 8'h1c;
			8'hc5: y = 8'ha6;
			8'hc6: y = 8'hb4;
			8'hc7: y = 8'hc6;
			8'hc8: y = 8'he8;
			8'hc9: y = 8'hdd;
			8'hca: y = 8'h74;
			8'hcb: y = 8'h1f;
			8'hcc: y = 8'h4b;
			8'hcd: y = 8'hbd;
			8'hce: y = 8'h8b;
			8'hcf: y = 8'h8a;
			8'hd0: y = 8'h70;
			8'hd1: y = 8'h3e;
			8'hd2: y = 8'hb5;
			8'hd3: y = 8'h66;
			8'hd4: y = 8'h48;
			8'hd5: y = 8'h03;
			8'hd6: y = 8'hf6;
			8'hd7: y = 8'h0e;
			8'hd8: y = 8'h61;
			8'hd9: y = 8'h35;
			8'hda: y = 8'h57;
			8'hdb: y = 8'hb9;
			8'hdc: y = 8'h86;
			8'hdd: y = 8'hc1;
			8'hde: y = 8'h1d;
			8'hdf: y = 8'h9e;
			8'he0: y = 8'he1;
			8'he1: y = 8'hf8;
			8'he2: y = 8'h98;
			8'he3: y = 8'h11;
			8'he4: y = 8'h69;
			8'he5: y = 8'hd9;
			8'he6: y = 8'h8e;
			8'he7: y = 8'h94;
			8'he8: y = 8'h9b;
			8'he9: y = 8'h1e;
			8'hea: y = 8'h87;
			8'heb: y = 8'he9;
			8'hec: y = 8'hce;
			8'hed: y = 8'h55;
			8'hee: y = 8'h28;
			8'hef: y = 8'hdf;
			8'hf0: y = 8'h8c;
			8'hf1: y = 8'ha1;
			8'hf2: y = 8'h89;
			8'hf3: y = 8'h0d;
			8'hf4: y = 8'hbf;
			8'hf5: y = 8'he6;
			8'hf6: y = 8'h42;
			8'hf7: y = 8'h68;
			8'hf8: y = 8'h41;
			8'hf9: y = 8'h99;
			8'hfa: y = 8'h2d;
			8'hfb: y = 8'h0f;
			8'hfc: y = 8'hb0;
			8'hfd: y = 8'h54;
			8'hfe: y = 8'hbb;
			8'hff: y = 8'h16;
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
module aesshiftrows64 (
	a,
	y
);
	input wire [127:0] a;
	output wire [63:0] y;
	assign y = {a[31:24], a[119:112], a[79:72], a[39:32], a[127:120], a[87:80], a[47:40], a[7:0]};
endmodule
module galoismultforward8 (
	a,
	y
);
	input wire [7:0] a;
	output wire [7:0] y;
	wire [7:0] leftshift;
	assign leftshift = {a[6:0], 1'b0};
	assign y = (a[7] ? leftshift ^ 8'b00011011 : leftshift);
endmodule
module galoismultinverse8 (
	a,
	y
);
	input wire [10:0] a;
	output wire [7:0] y;
	wire [7:0] temp0;
	wire [7:0] temp1;
	assign temp0 = (a[8] ? a[7:0] ^ 8'b00011011 : a[7:0]);
	assign temp1 = (a[9] ? temp0 ^ 8'b00110110 : temp0);
	assign y = (a[10] ? temp1 ^ 8'b01101100 : temp1);
endmodule
module rconlut32 (
	rd,
	rcon
);
	reg _sv2v_0;
	input wire [3:0] rd;
	output wire [31:0] rcon;
	reg [7:0] rcon8;
	always @(*) begin
		if (_sv2v_0)
			;
		case (rd)
			4'h0: rcon8 = 8'h01;
			4'h1: rcon8 = 8'h02;
			4'h2: rcon8 = 8'h04;
			4'h3: rcon8 = 8'h08;
			4'h4: rcon8 = 8'h10;
			4'h5: rcon8 = 8'h20;
			4'h6: rcon8 = 8'h40;
			4'h7: rcon8 = 8'h80;
			4'h8: rcon8 = 8'h1b;
			4'h9: rcon8 = 8'h36;
			4'ha: rcon8 = 8'h00;
			default: rcon8 = 8'h00;
		endcase
	end
	assign rcon = {24'b000000000000000000000000, rcon8};
	initial _sv2v_0 = 0;
endmodule
module rotate (
	a,
	shamt,
	y
);
	parameter WIDTH = 32;
	input wire [WIDTH - 1:0] a;
	input wire [$clog2(WIDTH) - 1:0] shamt;
	output wire [WIDTH - 1:0] y;
	assign y = (a << shamt) | (a >> (WIDTH - shamt));
endmodule
module bitmanipalu (
	A,
	B,
	W64,
	UW64,
	BSelect,
	ZBBSelect,
	Funct3,
	Funct7,
	Rs2E,
	LT,
	LTU,
	BALUControl,
	BMUActive,
	PreALUResult,
	FullResult,
	CondMaskB,
	CondShiftA,
	ALUResult
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[4216-:32]) - 1:0] A;
	input wire [$signed(P[4216-:32]) - 1:0] B;
	input wire W64;
	input wire UW64;
	input wire [3:0] BSelect;
	input wire [3:0] ZBBSelect;
	input wire [2:0] Funct3;
	input wire [6:0] Funct7;
	input wire [4:0] Rs2E;
	input wire LT;
	input wire LTU;
	input wire [2:0] BALUControl;
	input wire BMUActive;
	input wire [$signed(P[4216-:32]) - 1:0] PreALUResult;
	input wire [$signed(P[4216-:32]) - 1:0] FullResult;
	output wire [$signed(P[4216-:32]) - 1:0] CondMaskB;
	output wire [$signed(P[4216-:32]) - 1:0] CondShiftA;
	output reg [$signed(P[4216-:32]) - 1:0] ALUResult;
	wire [$signed(P[4216-:32]) - 1:0] ZBBResult;
	wire [$signed(P[4216-:32]) - 1:0] ZBCResult;
	wire [$signed(P[4216-:32]) - 1:0] ZBKBResult;
	wire [$signed(P[4216-:32]) - 1:0] ZBKXResult;
	wire [$signed(P[4216-:32]) - 1:0] ZKNHResult;
	wire [$signed(P[4216-:32]) - 1:0] ZKNDEResult;
	wire [$signed(P[4216-:32]) - 1:0] MaskB;
	wire [$signed(P[4216-:32]) - 1:0] RevA;
	wire Mask;
	wire PreShift;
	wire [1:0] PreShiftAmt;
	wire [$signed(P[4216-:32]) - 1:0] CondZextA;
	wire [$signed(P[4216-:32]) - 1:0] ABMU;
	wire [$signed(P[4216-:32]) - 1:0] BBMU;
	assign ABMU = A & {$signed(P[4216-:32]) {BMUActive}};
	assign BBMU = B & {$signed(P[4216-:32]) {BMUActive}};
	assign {Mask, PreShift} = BALUControl[1:0];
	generate
		if (P[1755]) begin : zbsdec
			decoder #(.BINARY_BITS($clog2($signed(P[4216-:32])))) maskgen(
				.binary(BBMU[$clog2($signed(P[4216-:32])) - 1:0]),
				.onehot(MaskB)
			);
			mux2 #(.WIDTH($signed(P[4216-:32]))) maskmux(
				.d0(B),
				.d1(MaskB),
				.s(Mask),
				.y(CondMaskB)
			);
		end
		else begin : genblk1
			assign CondMaskB = B;
		end
		if (P[1758]) begin : zbapreshift
			if ($signed(P[4216-:32]) == 64) begin : genblk1
				mux2 #(.WIDTH(64)) zextmux(
					.d0(A),
					.d1({{32 {1'b0}}, A[31:0]}),
					.s(UW64),
					.y(CondZextA)
				);
			end
			else begin : genblk1
				assign CondZextA = A;
			end
			assign PreShiftAmt = Funct3[2:1] & {2 {PreShift}};
			assign CondShiftA = CondZextA << PreShiftAmt;
		end
		else begin : genblk2
			assign PreShiftAmt = 2'b00;
			assign CondShiftA = A;
		end
		if ((P[1756] | P[1749]) | P[1757]) begin : bitreverse
			bitreverse #(.WIDTH($signed(P[4216-:32]))) brA(
				.A(ABMU),
				.RevA(RevA)
			);
		end
		if (P[1756] | P[1749]) begin : zbc
			zbc #(.P(P)) ZBC(
				.A(ABMU),
				.RevA(RevA),
				.B(BBMU),
				.Funct3(Funct3[1:0]),
				.ZBCResult(ZBCResult)
			);
		end
		else begin : genblk4
			assign ZBCResult = 1'sb0;
		end
		if (P[1757]) begin : zbb
			zbb #(.WIDTH($signed(P[4216-:32]))) ZBB(
				.A(ABMU),
				.RevA(RevA),
				.B(BBMU),
				.W64(W64),
				.LT(LT),
				.LTU(LTU),
				.BUnsigned(Funct3[0]),
				.ZBBSelect(ZBBSelect[2:0]),
				.ZBBResult(ZBBResult)
			);
		end
		else if (P[1750]) begin : zbkbonly
			genvar _gv_i_8;
			for (_gv_i_8 = 0; _gv_i_8 < $signed(P[4216-:32]); _gv_i_8 = _gv_i_8 + 8) begin : byteloop
				localparam i = _gv_i_8;
				assign ZBBResult[($signed(P[4216-:32]) - i) - 1:($signed(P[4216-:32]) - i) - 8] = ABMU[i + 7:i];
			end
		end
		else begin : genblk5
			assign ZBBResult = 1'sb0;
		end
		if (P[1750]) begin : zbkb
			zbkb #(.WIDTH($signed(P[4216-:32]))) ZBKB(
				.A(ABMU),
				.B(BBMU[($signed(P[4216-:32]) / 2) - 1:0]),
				.Funct3(Funct3),
				.ZBKBSelect(ZBBSelect[2:0]),
				.ZBKBResult(ZBKBResult)
			);
		end
		else begin : genblk6
			assign ZBKBResult = 1'sb0;
		end
		if (P[1748]) begin : zbkx
			zbkx #(.WIDTH($signed(P[4216-:32]))) ZBKX(
				.A(ABMU),
				.B(BBMU),
				.ZBKXSelect(ZBBSelect[0]),
				.ZBKXResult(ZBKXResult)
			);
		end
		else begin : genblk7
			assign ZBKXResult = 1'sb0;
		end
		if (P[1747] | P[1746]) begin : zknde
			if ($signed(P[4216-:32]) == 32) begin : genblk1
				zknde32 #(.P(P)) ZKN32(
					.A(ABMU),
					.B(BBMU),
					.bs(Funct7[6:5]),
					.round(Rs2E[3:0]),
					.ZKNSelect(ZBBSelect[3:0]),
					.ZKNDEResult(ZKNDEResult)
				);
			end
			else begin : genblk1
				zknde64 #(.P(P)) ZKN64(
					.A(ABMU),
					.B(BBMU),
					.round(Rs2E[3:0]),
					.ZKNSelect(ZBBSelect[3:0]),
					.ZKNDEResult(ZKNDEResult)
				);
			end
		end
		else begin : genblk8
			assign ZKNDEResult = 1'sb0;
		end
		if (P[1745]) begin : zknh
			if ($signed(P[4216-:32]) == 32) begin : genblk1
				zknh32 ZKNH32(
					.A(ABMU),
					.B(BBMU),
					.ZKNHSelect(ZBBSelect),
					.ZKNHResult(ZKNHResult)
				);
			end
			else begin : genblk1
				zknh64 ZKNH64(
					.A(ABMU),
					.ZKNHSelect(ZBBSelect),
					.ZKNHResult(ZKNHResult)
				);
			end
		end
		else begin : genblk9
			assign ZKNHResult = 1'sb0;
		end
	endgenerate
	always @(*) begin
		if (_sv2v_0)
			;
		case (BSelect)
			4'b0000: ALUResult = PreALUResult;
			4'b0001: ALUResult = FullResult;
			4'b0010: ALUResult = ZBBResult;
			4'b0011: ALUResult = ZBCResult;
			4'b0100: ALUResult = ZBKBResult;
			4'b0110: ALUResult = ZBKXResult;
			4'b0111: ALUResult = ZKNDEResult;
			4'b1000: ALUResult = ZKNHResult;
			default: ALUResult = PreALUResult;
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
module bitreverse (
	A,
	RevA
);
	parameter WIDTH = 32;
	input wire [WIDTH - 1:0] A;
	output wire [WIDTH - 1:0] RevA;
	genvar _gv_i_9;
	generate
		for (_gv_i_9 = 0; _gv_i_9 < WIDTH; _gv_i_9 = _gv_i_9 + 1) begin : loop
			localparam i = _gv_i_9;
			assign RevA[(WIDTH - i) - 1] = A[i];
		end
	endgenerate
endmodule
module bmuctrl (
	clk,
	reset,
	InstrD,
	ALUOpD,
	BRegWriteD,
	BALUSrcBD,
	BW64D,
	BUW64D,
	BSubArithD,
	IllegalBitmanipInstrD,
	StallE,
	FlushE,
	ALUSelectD,
	BSelectE,
	ZBBSelectE,
	BALUControlE,
	BMUActiveE
);
	reg _sv2v_0;
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire [31:0] InstrD;
	input wire ALUOpD;
	output wire BRegWriteD;
	output wire BALUSrcBD;
	output wire BW64D;
	output wire BUW64D;
	output wire BSubArithD;
	output wire IllegalBitmanipInstrD;
	input wire StallE;
	input wire FlushE;
	output wire [2:0] ALUSelectD;
	output wire [3:0] BSelectE;
	output wire [3:0] ZBBSelectE;
	output wire [2:0] BALUControlE;
	output wire BMUActiveE;
	wire [6:0] OpD;
	wire [2:0] Funct3D;
	wire [6:0] Funct7D;
	wire [4:0] Rs2D;
	wire RotateD;
	wire MaskD;
	wire PreShiftD;
	wire [2:0] BALUControlD;
	wire [2:0] BALUSelectD;
	wire BALUOpD;
	wire [3:0] BSelectD;
	wire [3:0] ZBBSelectD;
	reg [20:0] BMUControlsD;
	assign OpD = InstrD[6:0];
	assign Funct3D = InstrD[14:12];
	assign Funct7D = InstrD[31:25];
	assign Rs2D = InstrD[24:20];
	always @(*) begin
		if (_sv2v_0)
			;
		BMUControlsD = 21'b000000000000000000001;
		if (P[1758]) begin
			casez ({OpD, Funct7D, Funct3D})
				17'b01100110010000010: BMUControlsD = 21'b000000100001000100010;
				17'b01100110010000100: BMUControlsD = 21'b000000100001000100010;
				17'b01100110010000110: BMUControlsD = 21'b000000100001000100010;
			endcase
			if ($signed(P[4216-:32]) == 64)
				casez ({OpD, Funct7D, Funct3D})
					17'b01110110010000010: BMUControlsD = 21'b000000100001001100010;
					17'b01110110010000100: BMUControlsD = 21'b000000100001001100010;
					17'b01110110010000110: BMUControlsD = 21'b000000100001001100010;
					17'b01110110000100000: BMUControlsD = 21'b000000100001001100000;
					17'b0011011000010z001: BMUControlsD = 21'b001000100001101100000;
				endcase
		end
		if (P[1757]) begin
			casez ({OpD, Funct7D, Funct3D})
				17'b00100110110000001:
					if (Rs2D[4:1] == 4'b0010)
						BMUControlsD = 21'b000001000011100100000;
					else if ((Rs2D[4:2] == 3'b000) & ~(Rs2D[1] & Rs2D[0]))
						BMUControlsD = 21'b000001000001100100000;
				17'b00100110010100101:
					if (Rs2D[4:0] == 5'b00111)
						BMUControlsD = 21'b000001000101100100000;
				17'b01100110000101110: BMUControlsD = 21'b000001001111000110000;
				17'b01100110000101111: BMUControlsD = 21'b000001001111000110000;
				17'b01100110000101100: BMUControlsD = 21'b000001000111000110000;
				17'b01100110000101101: BMUControlsD = 21'b000001000111000110000;
			endcase
			if ($signed(P[4216-:32]) == 32)
				casez ({OpD, Funct7D, Funct3D})
					17'b01100110000100100: BMUControlsD = 21'b000001000011100100000;
				endcase
			else if ($signed(P[4216-:32]) == 64)
				casez ({OpD, Funct7D, Funct3D})
					17'b01110110000100100: BMUControlsD = 21'b000001000011000100000;
					17'b00110110110000001:
						if ((Rs2D[4:2] == 3'b000) & ~(Rs2D[1] & Rs2D[0]))
							BMUControlsD = 21'b000001000001111000000;
				endcase
		end
		if (P[1756])
			casez ({OpD, Funct7D, Funct3D})
				17'b01100110000101010: BMUControlsD = 21'b000001100011000100000;
				17'b011001100001010z1: BMUControlsD = 21'b000001100001000100000;
			endcase
		if (P[1749])
			casez ({OpD, Funct7D, Funct3D})
				17'b011001100001010z1: BMUControlsD = 21'b000001100001000100000;
			endcase
		if (P[1755]) begin
			casez ({OpD, Funct7D, Funct3D})
				17'b01100110100100001: BMUControlsD = 21'b111000100001000110100;
				17'b01100110100100101: BMUControlsD = 21'b101000100001000100100;
				17'b01100110110100001: BMUControlsD = 21'b100000100001000100100;
				17'b01100110010100001: BMUControlsD = 21'b110000100001000100100;
			endcase
			if ($signed(P[4216-:32]) == 32)
				casez ({OpD, Funct7D, Funct3D})
					17'b00100110100100001: BMUControlsD = 21'b111000100001100110100;
					17'b00100110100100101: BMUControlsD = 21'b101000100001100100100;
					17'b00100110110100001: BMUControlsD = 21'b100000100001100100100;
					17'b00100110010100001: BMUControlsD = 21'b110000100001100100100;
				endcase
			else if ($signed(P[4216-:32]) == 64)
				casez ({OpD, Funct7D, Funct3D})
					17'b0010011010010z001: BMUControlsD = 21'b111000100001100110100;
					17'b0010011010010z101: BMUControlsD = 21'b101000100001100100100;
					17'b0010011011010z001: BMUControlsD = 21'b100000100001100100100;
					17'b0010011001010z001: BMUControlsD = 21'b110000100001100100100;
				endcase
		end
		if (P[1757] | P[1755])
			casez ({OpD, Funct7D, Funct3D})
				17'b01100110000000001: BMUControlsD = 21'b001000000001000100000;
				17'b01100110z00000101: BMUControlsD = 21'b001000000001000100000;
				17'b0010011000000z001:
					if (($signed(P[4216-:32]) == 64) | !Funct7D[0])
						BMUControlsD = 21'b001000000001100100000;
				17'b00100110z0000z101:
					if (($signed(P[4216-:32]) == 64) | !Funct7D[0])
						BMUControlsD = 21'b001000000001100100000;
				17'b01110110000000001:
					if ($signed(P[4216-:32]) == 64)
						BMUControlsD = 21'b001000000001010100000;
				17'b01110110z00000101:
					if ($signed(P[4216-:32]) == 64)
						BMUControlsD = 21'b001000000001010100000;
				17'b00110110000000001:
					if ($signed(P[4216-:32]) == 64)
						BMUControlsD = 21'b001000000001110100000;
				17'b00110110z00000101:
					if ($signed(P[4216-:32]) == 64)
						BMUControlsD = 21'b001000000001110100000;
			endcase
		if (P[1750]) begin
			casez ({OpD, Funct7D, Funct3D})
				17'b01100110000100100: BMUControlsD = 21'b000010000011000100000;
				17'b01100110000100111: BMUControlsD = 21'b000010000011000100000;
				17'b00100110110100101:
					if (Rs2D == 5'b00111)
						BMUControlsD = 21'b000010000001100100000;
			endcase
			if ($signed(P[4216-:32]) == 32)
				casez ({OpD, Funct7D, Funct3D})
					17'b00100110000100001:
						if (Rs2D == 5'b01111)
							BMUControlsD = 21'b000010000111100100000;
					17'b00100110000100101:
						if (Rs2D == 5'b01111)
							BMUControlsD = 21'b000010000111100100000;
				endcase
			else if ($signed(P[4216-:32]) == 64)
				casez ({OpD, Funct7D, Funct3D})
					17'b01110110000100100: BMUControlsD = 21'b000010001011010100000;
				endcase
		end
		if (P[1757] | P[1750]) begin
			casez ({OpD, Funct7D, Funct3D})
				17'b01100110110000001: BMUControlsD = 21'b001000101111000101000;
				17'b01100110110000101: BMUControlsD = 21'b001000101111000101000;
				17'b01100110100000111: BMUControlsD = 21'b111000101111000110000;
				17'b01100110100000110: BMUControlsD = 21'b110000101111000110000;
				17'b01100110100000100: BMUControlsD = 21'b100000101111000110000;
				17'b0010011011010z101:
					if ((($signed(P[4216-:32]) == 32) ^ Funct7D[0]) & (Rs2D == 5'b11000))
						BMUControlsD = 21'b000001000101100100000;
			endcase
			if ($signed(P[4216-:32]) == 32)
				casez ({OpD, Funct7D, Funct3D})
					17'b00100110110000101: BMUControlsD = 21'b001000001111100101000;
				endcase
			else if ($signed(P[4216-:32]) == 64)
				casez ({OpD, Funct7D, Funct3D})
					17'b01110110110000001: BMUControlsD = 21'b001000001111010101000;
					17'b01110110110000101: BMUControlsD = 21'b001000001111010101000;
					17'b0010011011000z101: BMUControlsD = 21'b001000001111100101000;
					17'b00110110110000101: BMUControlsD = 21'b001000001111110101000;
				endcase
		end
		if (P[1748])
			casez ({OpD, Funct7D, Funct3D})
				17'b01100110010100100: BMUControlsD = 21'b000011000001000100000;
				17'b01100110010100010: BMUControlsD = 21'b000011000011000100000;
			endcase
		if (P[1747]) begin
			if ($signed(P[4216-:32]) == 32)
				casez ({OpD, Funct7D, Funct3D})
					17'b0110011zz10101000: BMUControlsD = 21'b000011101001000100000;
					17'b0110011zz10111000: BMUControlsD = 21'b000011100001000100000;
				endcase
			else if ($signed(P[4216-:32]) == 64)
				casez ({OpD, Funct7D, Funct3D})
					17'b01100110011101000: BMUControlsD = 21'b000011101001000100000;
					17'b01100110011111000: BMUControlsD = 21'b000011100001000100000;
					17'b00100110011000001:
						if (Rs2D == 5'b00000)
							BMUControlsD = 21'b000011110001100100000;
				endcase
		end
		if (P[1746]) begin
			if ($signed(P[4216-:32]) == 32)
				casez ({OpD, Funct7D, Funct3D})
					17'b0110011zz10001000: BMUControlsD = 21'b000011101011000100000;
					17'b0110011zz10011000: BMUControlsD = 21'b000011100011000100000;
				endcase
			else if ($signed(P[4216-:32]) == 64)
				casez ({OpD, Funct7D, Funct3D})
					17'b01100110011001000: BMUControlsD = 21'b000011101011000100000;
					17'b01100110011011000: BMUControlsD = 21'b000011100011000100000;
				endcase
		end
		if ((P[1747] | P[1746]) & ($signed(P[4216-:32]) == 64))
			casez ({OpD, Funct7D, Funct3D})
				17'b00100110011000001:
					if ((Rs2D[4] == 1'b1) & ($unsigned(Rs2D[3:0]) <= 10))
						BMUControlsD = 21'b000011100101000100000;
				17'b01100110111111000: BMUControlsD = 21'b000011100111000100000;
			endcase
		if (P[1745]) begin
			casez ({OpD, Funct7D, Funct3D})
				17'b00100110001000001:
					if (Rs2D == 5'b00010)
						BMUControlsD = 21'b000100000001000100000;
					else if (Rs2D == 5'b00011)
						BMUControlsD = 21'b000100000011000100000;
					else if (Rs2D == 5'b00000)
						BMUControlsD = 21'b000100000101000100000;
					else if (Rs2D == 5'b00001)
						BMUControlsD = 21'b000100000111000100000;
			endcase
			if ($signed(P[4216-:32]) == 32)
				casez ({OpD, Funct7D, Funct3D})
					17'b01100110101110000: BMUControlsD = 21'b000100010001000100000;
					17'b01100110101010000: BMUControlsD = 21'b000100010011000100000;
					17'b01100110101111000: BMUControlsD = 21'b000100010101000100000;
					17'b01100110101011000: BMUControlsD = 21'b000100010111000100000;
					17'b01100110101000000: BMUControlsD = 21'b000100011001000100000;
					17'b01100110101001000: BMUControlsD = 21'b000100011101000100000;
				endcase
			else if ($signed(P[4216-:32]) == 64)
				casez ({OpD, Funct7D, Funct3D})
					17'b00100110001000001:
						if (Rs2D == 5'b00110)
							BMUControlsD = 21'b000100010001000100000;
						else if (Rs2D == 5'b00111)
							BMUControlsD = 21'b000100010011000100000;
						else if (Rs2D == 5'b00100)
							BMUControlsD = 21'b000100010101000100000;
						else if (Rs2D == 5'b00101)
							BMUControlsD = 21'b000100010111000100000;
				endcase
		end
	end
	assign {BALUSelectD, BSelectD, ZBBSelectD, BRegWriteD, BALUSrcBD, BW64D, BUW64D, BALUOpD, BSubArithD, RotateD, MaskD, PreShiftD, IllegalBitmanipInstrD} = BMUControlsD;
	assign BALUControlD = {RotateD, MaskD, PreShiftD};
	assign ALUSelectD = (BALUOpD ? BALUSelectD : (ALUOpD ? Funct3D : 3'b000));
	flopenrc #(.WIDTH(12)) controlregBMU(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d({BSelectD, ZBBSelectD, BALUControlD, ~IllegalBitmanipInstrD}),
		.q({BSelectE, ZBBSelectE, BALUControlE, BMUActiveE})
	);
	initial _sv2v_0 = 0;
endmodule
module byteop (
	A,
	ByteSelect,
	ByteResult
);
	parameter WIDTH = 32;
	input wire [WIDTH - 1:0] A;
	input wire ByteSelect;
	output wire [WIDTH - 1:0] ByteResult;
	wire [WIDTH - 1:0] OrcBResult;
	wire [WIDTH - 1:0] Rev8Result;
	genvar _gv_i_10;
	generate
		for (_gv_i_10 = 0; _gv_i_10 < WIDTH; _gv_i_10 = _gv_i_10 + 8) begin : byteloop
			localparam i = _gv_i_10;
			assign OrcBResult[i + 7:i] = {8 {|A[i + 7:i]}};
			assign Rev8Result[(WIDTH - i) - 1:(WIDTH - i) - 8] = A[i + 7:i];
		end
	endgenerate
	mux2 #(.WIDTH(WIDTH)) byteresultmux(
		.d0(Rev8Result),
		.d1(OrcBResult),
		.s(ByteSelect),
		.y(ByteResult)
	);
endmodule
module clmul (
	X,
	Y,
	ClmulResult
);
	reg _sv2v_0;
	parameter WIDTH = 32;
	input wire [WIDTH - 1:0] X;
	input wire [WIDTH - 1:0] Y;
	output reg [WIDTH - 1:0] ClmulResult;
	reg [(WIDTH * WIDTH) - 1:0] S;
	integer i;
	integer j;
	always @(*) begin
		if (_sv2v_0)
			;
		for (i = 0; i < WIDTH; i = i + 1)
			begin : outer
				S[WIDTH * i] = X[0] & Y[i];
				for (j = 1; j <= i; j = j + 1)
					begin : inner
						S[(WIDTH * i) + j] = (X[j] & Y[i - j]) ^ S[((WIDTH * i) + j) - 1];
					end
				ClmulResult[i] = S[((WIDTH * i) + j) - 1];
			end
	end
	initial _sv2v_0 = 0;
endmodule
module cnt (
	A,
	RevA,
	B,
	W64,
	CntResult
);
	parameter WIDTH = 32;
	input wire [WIDTH - 1:0] A;
	input wire [WIDTH - 1:0] RevA;
	input wire [1:0] B;
	input wire W64;
	output wire [WIDTH - 1:0] CntResult;
	wire [WIDTH - 1:0] czResult;
	wire [WIDTH - 1:0] cpopResult;
	wire [WIDTH - 1:0] lzcA;
	wire [WIDTH - 1:0] popcntA;
	generate
		if (WIDTH == 64) begin : genblk1
			mux4 #(.WIDTH(WIDTH)) lzcmux64(
				.d0(A),
				.d1({A[31:0], {32 {1'b1}}}),
				.d2(RevA),
				.d3({RevA[63:32], {32 {1'b1}}}),
				.s({B[0], W64}),
				.y(lzcA)
			);
			mux2 #(.WIDTH(WIDTH)) popcntmux64(
				.d0(A),
				.d1({{32 {1'b0}}, A[31:0]}),
				.s(W64),
				.y(popcntA)
			);
		end
		else begin : genblk1
			assign popcntA = A;
			mux2 #(.WIDTH(WIDTH)) lzcmux32(
				.d0(A),
				.d1(RevA),
				.s(B[0]),
				.y(lzcA)
			);
		end
	endgenerate
	lzc #(.WIDTH(WIDTH)) lzc(
		.num(lzcA),
		.ZeroCnt(czResult[$clog2(WIDTH):0])
	);
	popcnt #(.WIDTH(WIDTH)) popcntw(
		.num(popcntA),
		.PopCnt(cpopResult[$clog2(WIDTH):0])
	);
	assign czResult[WIDTH - 1:$clog2(WIDTH) + 1] = 1'sb0;
	assign cpopResult[WIDTH - 1:$clog2(WIDTH) + 1] = 1'sb0;
	mux2 #(.WIDTH(WIDTH)) cntresultmux(
		.d0(czResult),
		.d1(cpopResult),
		.s(B[1]),
		.y(CntResult)
	);
endmodule
module ext (
	A,
	ExtSelect,
	ExtResult
);
	parameter WIDTH = 32;
	input wire [15:0] A;
	input wire [1:0] ExtSelect;
	output wire [WIDTH - 1:0] ExtResult;
	wire [WIDTH - 1:0] sexthResult;
	wire [WIDTH - 1:0] zexthResult;
	wire [WIDTH - 1:0] sextbResult;
	assign sexthResult = {{WIDTH - 16 {A[15]}}, A[15:0]};
	assign zexthResult = {{WIDTH - 16 {1'b0}}, A[15:0]};
	assign sextbResult = {{WIDTH - 8 {A[7]}}, A[7:0]};
	mux3 #(.WIDTH(WIDTH)) extmux(
		.d0(sextbResult),
		.d1(sexthResult),
		.d2(zexthResult),
		.s(ExtSelect),
		.y(ExtResult)
	);
endmodule
module popcnt (
	num,
	PopCnt
);
	reg _sv2v_0;
	parameter WIDTH = 32;
	input wire [WIDTH - 1:0] num;
	output wire [$clog2(WIDTH):0] PopCnt;
	reg [$clog2(WIDTH):0] sum;
	always @(*) begin
		if (_sv2v_0)
			;
		sum = 1'sb0;
		begin : sv2v_autoblock_1
			reg signed [31:0] i;
			for (i = 0; i < WIDTH; i = i + 1)
				begin : loop
					sum = (num[i] ? sum + 1 : sum);
				end
		end
	end
	assign PopCnt = sum;
	initial _sv2v_0 = 0;
endmodule
module zbb (
	A,
	RevA,
	B,
	W64,
	LT,
	LTU,
	BUnsigned,
	ZBBSelect,
	ZBBResult
);
	parameter WIDTH = 32;
	input wire [WIDTH - 1:0] A;
	input wire [WIDTH - 1:0] RevA;
	input wire [WIDTH - 1:0] B;
	input wire W64;
	input wire LT;
	input wire LTU;
	input wire BUnsigned;
	input wire [2:0] ZBBSelect;
	output wire [WIDTH - 1:0] ZBBResult;
	wire lt;
	wire [WIDTH - 1:0] CntResult;
	wire [WIDTH - 1:0] MinMaxResult;
	wire [WIDTH - 1:0] ByteResult;
	wire [WIDTH - 1:0] ExtResult;
	mux2 #(.WIDTH(1)) ltmux(
		.d0(LT),
		.d1(LTU),
		.s(BUnsigned),
		.y(lt)
	);
	cnt #(.WIDTH(WIDTH)) cnt(
		.A(A),
		.RevA(RevA),
		.B(B[1:0]),
		.W64(W64),
		.CntResult(CntResult)
	);
	byteop #(.WIDTH(WIDTH)) bu(
		.A(A),
		.ByteSelect(B[0]),
		.ByteResult(ByteResult)
	);
	ext #(.WIDTH(WIDTH)) ext(
		.A(A[15:0]),
		.ExtSelect({~B[2], B[2] & B[0]}),
		.ExtResult(ExtResult)
	);
	mux2 #(.WIDTH(WIDTH)) minmaxmux(
		.d0(B),
		.d1(A),
		.s(ZBBSelect[2] ^ lt),
		.y(MinMaxResult)
	);
	mux4 #(.WIDTH(WIDTH)) zbbresultmux(
		.d0(CntResult),
		.d1(ExtResult),
		.d2(ByteResult),
		.d3(MinMaxResult),
		.s(ZBBSelect[1:0]),
		.y(ZBBResult)
	);
endmodule
module zbc (
	A,
	RevA,
	B,
	Funct3,
	ZBCResult
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[4216-:32]) - 1:0] A;
	input wire [$signed(P[4216-:32]) - 1:0] RevA;
	input wire [$signed(P[4216-:32]) - 1:0] B;
	input wire [1:0] Funct3;
	output wire [$signed(P[4216-:32]) - 1:0] ZBCResult;
	wire [$signed(P[4216-:32]) - 1:0] ClmulResult;
	wire [$signed(P[4216-:32]) - 1:0] RevClmulResult;
	wire [$signed(P[4216-:32]) - 1:0] RevB;
	wire [$signed(P[4216-:32]) - 1:0] X;
	wire [$signed(P[4216-:32]) - 1:0] Y;
	bitreverse #(.WIDTH($signed(P[4216-:32]))) brB(
		.A(B),
		.RevA(RevB)
	);
	generate
		if (P[1756]) begin : genblk1
			mux3 #(.WIDTH($signed(P[4216-:32]))) xmux(
				.d0({RevA[$signed(P[4216-:32]) - 2:0], 1'b0}),
				.d1(RevA),
				.d2(A),
				.s(~Funct3[1:0]),
				.y(X)
			);
		end
		else begin : genblk1
			mux2 #(.WIDTH($signed(P[4216-:32]))) xmux(
				.d0(A),
				.d1({RevA[$signed(P[4216-:32]) - 2:0], 1'b0}),
				.s(Funct3[1]),
				.y(X)
			);
		end
	endgenerate
	mux2 #(.WIDTH($signed(P[4216-:32]))) ymux(
		.d0(B),
		.d1(RevB),
		.s(Funct3[1]),
		.y(Y)
	);
	clmul #(.WIDTH($signed(P[4216-:32]))) clm(
		.X(X),
		.Y(Y),
		.ClmulResult(ClmulResult)
	);
	bitreverse #(.WIDTH($signed(P[4216-:32]))) brClmulResult(
		.A(ClmulResult),
		.RevA(RevClmulResult)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) zbcresultmux(
		.d0(ClmulResult),
		.d1(RevClmulResult),
		.s(Funct3[1]),
		.y(ZBCResult)
	);
endmodule
module packer (
	A,
	B,
	PackSelect,
	PackResult
);
	reg _sv2v_0;
	parameter WIDTH = 32;
	input wire [(WIDTH / 2) - 1:0] A;
	input wire [(WIDTH / 2) - 1:0] B;
	input wire [2:0] PackSelect;
	output reg [WIDTH - 1:0] PackResult;
	wire [(WIDTH / 2) - 1:0] lowhalf;
	wire [(WIDTH / 2) - 1:0] highhalf;
	wire [7:0] lowhalfh;
	wire [7:0] highhalfh;
	wire [15:0] lowhalfw;
	wire [15:0] highhalfw;
	wire [WIDTH - 1:0] Pack;
	wire [WIDTH - 1:0] PackH;
	wire [WIDTH - 1:0] PackW;
	assign lowhalf = A[(WIDTH / 2) - 1:0];
	assign highhalf = B[(WIDTH / 2) - 1:0];
	assign lowhalfh = A[7:0];
	assign highhalfh = B[7:0];
	assign lowhalfw = A[15:0];
	assign highhalfw = B[15:0];
	assign Pack = {highhalf, lowhalf};
	assign PackH = {{WIDTH - 16 {1'b0}}, highhalfh, lowhalfh};
	assign PackW = (WIDTH == 64 ? {{WIDTH - 32 {highhalfw[15]}}, highhalfw, lowhalfw} : Pack);
	always @(*) begin
		if (_sv2v_0)
			;
		if (PackSelect[1:0] == 2'b11)
			PackResult = PackH;
		else if (PackSelect[2] == 1'b0)
			PackResult = Pack;
		else
			PackResult = PackW;
	end
	initial _sv2v_0 = 0;
endmodule
module zbkb (
	A,
	B,
	Funct3,
	ZBKBSelect,
	ZBKBResult
);
	parameter WIDTH = 32;
	input wire [WIDTH - 1:0] A;
	input wire [(WIDTH / 2) - 1:0] B;
	input wire [2:0] Funct3;
	input wire [2:0] ZBKBSelect;
	output wire [WIDTH - 1:0] ZBKBResult;
	wire [WIDTH - 1:0] Brev8Result;
	wire [WIDTH - 1:0] PackResult;
	wire [WIDTH - 1:0] ZipResult;
	genvar _gv_i_11;
	genvar _gv_j_1;
	generate
		for (_gv_i_11 = 0; _gv_i_11 < (WIDTH / 8); _gv_i_11 = _gv_i_11 + 1) begin : genblk1
			localparam i = _gv_i_11;
			for (_gv_j_1 = 0; _gv_j_1 < 8; _gv_j_1 = _gv_j_1 + 1) begin : genblk1
				localparam j = _gv_j_1;
				assign Brev8Result[(i * 8) + j] = A[((i * 8) + 7) - j];
			end
		end
	endgenerate
	packer #(.WIDTH(WIDTH)) pack(
		.A(A[(WIDTH / 2) - 1:0]),
		.B(B[(WIDTH / 2) - 1:0]),
		.PackSelect({ZBKBSelect[2], Funct3[1:0]}),
		.PackResult(PackResult)
	);
	zipper #(.WIDTH(WIDTH)) zipper(
		.A(A),
		.ZipSelect(Funct3[2]),
		.ZipResult(ZipResult)
	);
	mux3 #(.WIDTH(WIDTH)) zbkbresultmux(
		.d0(Brev8Result),
		.d1(PackResult),
		.d2(ZipResult),
		.s(ZBKBSelect[1:0]),
		.y(ZBKBResult)
	);
endmodule
module zbkx (
	A,
	B,
	ZBKXSelect,
	ZBKXResult
);
	reg _sv2v_0;
	parameter WIDTH = 32;
	input wire [WIDTH - 1:0] A;
	input wire [WIDTH - 1:0] B;
	input wire ZBKXSelect;
	output wire [WIDTH - 1:0] ZBKXResult;
	reg [WIDTH - 1:0] xperm4;
	reg [WIDTH - 1:0] xperm8;
	reg [WIDTH - 1:0] xperm4lookup;
	reg [WIDTH - 1:0] xperm8lookup;
	reg signed [31:0] i;
	always @(*) begin
		if (_sv2v_0)
			;
		for (i = 0; i < WIDTH; i = i + 4)
			begin : xperm4calc
				xperm4lookup = A >> {B[i+:4], 2'b00};
				xperm4[i+:4] = xperm4lookup[3:0];
			end
		for (i = 0; i < WIDTH; i = i + 8)
			begin : xperm8calc
				xperm8lookup = A >> {B[i+:8], 3'b000};
				xperm8[i+:8] = xperm8lookup[7:0];
			end
	end
	assign ZBKXResult = (ZBKXSelect ? xperm4 : xperm8);
	initial _sv2v_0 = 0;
endmodule
module zipper (
	A,
	ZipSelect,
	ZipResult
);
	parameter WIDTH = 64;
	input wire [WIDTH - 1:0] A;
	input wire ZipSelect;
	output wire [WIDTH - 1:0] ZipResult;
	wire [WIDTH - 1:0] zip;
	wire [WIDTH - 1:0] unzip;
	genvar _gv_i_12;
	generate
		for (_gv_i_12 = 0; _gv_i_12 < (WIDTH / 2); _gv_i_12 = _gv_i_12 + 1) begin : loop
			localparam i = _gv_i_12;
			assign zip[2 * i] = A[i];
			assign zip[(2 * i) + 1] = A[i + (WIDTH / 2)];
			assign unzip[i] = A[2 * i];
			assign unzip[i + (WIDTH / 2)] = A[(2 * i) + 1];
		end
	endgenerate
	mux2 #(.WIDTH(WIDTH)) ZipMux(
		.d0(zip),
		.d1(unzip),
		.s(ZipSelect),
		.y(ZipResult)
	);
endmodule
module zknde32 (
	A,
	B,
	bs,
	round,
	ZKNSelect,
	ZKNDEResult
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [31:0] A;
	input wire [31:0] B;
	input wire [1:0] bs;
	input wire [3:0] round;
	input wire [3:0] ZKNSelect;
	output wire [31:0] ZKNDEResult;
	wire [4:0] shamt;
	wire [7:0] SboxIn;
	wire [31:0] ZKNEResult;
	wire [31:0] ZKNDResult;
	wire [31:0] rotin;
	wire [31:0] rotout;
	assign shamt = {bs, 3'b000};
	assign SboxIn = B[shamt+:8];
	generate
		if (P[1747]) begin : genblk1
			aes32d aes32d(
				.SboxIn(SboxIn),
				.finalround(ZKNSelect[2]),
				.result(ZKNDResult)
			);
		end
		if (P[1746]) begin : genblk2
			aes32e aes32e(
				.SboxIn(SboxIn),
				.finalround(ZKNSelect[2]),
				.result(ZKNEResult)
			);
		end
		if (P[1747] & P[1746]) begin : genblk3
			mux2 #(.WIDTH(32)) zknmux(
				.d0(ZKNDResult),
				.d1(ZKNEResult),
				.s(ZKNSelect[0]),
				.y(rotin)
			);
		end
		else if (P[1747]) begin : genblk3
			assign rotin = ZKNDResult;
		end
		else begin : genblk3
			assign rotin = ZKNEResult;
		end
	endgenerate
	mux4 #(.WIDTH(32)) mrotmux(
		.d0(rotin),
		.d1({rotin[23:0], rotin[31:24]}),
		.d2({rotin[15:0], rotin[31:16]}),
		.d3({rotin[7:0], rotin[31:8]}),
		.s(bs),
		.y(rotout)
	);
	assign ZKNDEResult = A ^ rotout;
endmodule
module zknde64 (
	A,
	B,
	round,
	ZKNSelect,
	ZKNDEResult
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [63:0] A;
	input wire [63:0] B;
	input wire [3:0] round;
	input wire [3:0] ZKNSelect;
	output wire [63:0] ZKNDEResult;
	wire [63:0] aes64dRes;
	wire [63:0] aes64eRes;
	wire [63:0] aes64ks1iRes;
	wire [63:0] aes64ks2Res;
	wire [31:0] SboxEIn;
	wire [31:0] SboxKIn;
	wire [31:0] Sbox0In;
	wire [31:0] Sbox0Out;
	generate
		if (P[1747]) begin : genblk1
			aes64d aes64d(
				.rs1(A),
				.rs2(B),
				.finalround(ZKNSelect[2]),
				.aes64im(ZKNSelect[3]),
				.result(aes64dRes)
			);
		end
		else begin : genblk1
			assign aes64dRes = 1'sb0;
		end
		if (P[1746]) begin : genblk2
			aes64e aes64e(
				.rs1(A),
				.rs2(B),
				.finalround(ZKNSelect[2]),
				.Sbox0Out(Sbox0Out),
				.SboxEIn(SboxEIn),
				.result(aes64eRes)
			);
			mux2 #(.WIDTH(32)) sboxmux(
				.d0(SboxEIn),
				.d1(SboxKIn),
				.s(ZKNSelect[1]),
				.y(Sbox0In)
			);
		end
		else begin : genblk2
			assign aes64eRes = 1'sb0;
			assign Sbox0In = SboxKIn;
		end
	endgenerate
	aessbox32 sbox(
		.a(Sbox0In),
		.y(Sbox0Out)
	);
	aes64ks1i aes64ks1i(
		.round(round),
		.rs1(A[63:32]),
		.Sbox0Out(Sbox0Out),
		.SboxKIn(SboxKIn),
		.result(aes64ks1iRes)
	);
	aes64ks2 aes64ks2(
		.rs2(B),
		.rs1(A[63:32]),
		.result(aes64ks2Res)
	);
	mux4 #(.WIDTH(64)) zkndmux(
		.d0(aes64dRes),
		.d1(aes64eRes),
		.d2(aes64ks1iRes),
		.d3(aes64ks2Res),
		.s(ZKNSelect[1:0]),
		.y(ZKNDEResult)
	);
endmodule
module zknh32 (
	A,
	B,
	ZKNHSelect,
	ZKNHResult
);
	input wire [31:0] A;
	input wire [31:0] B;
	input wire [3:0] ZKNHSelect;
	output wire [31:0] ZKNHResult;
	wire [31:0] sha256res;
	wire [31:0] sha512res;
	sha256 sha256(
		.A(A),
		.ZKNHSelect(ZKNHSelect[1:0]),
		.result(sha256res)
	);
	sha512_32 sha512(
		.A(A),
		.B(B),
		.ZKNHSelect(ZKNHSelect[2:0]),
		.result(sha512res)
	);
	mux2 #(.WIDTH(32)) resultmux(
		.d0(sha256res),
		.d1(sha512res),
		.s(ZKNHSelect[3]),
		.y(ZKNHResult)
	);
endmodule
module zknh64 (
	A,
	ZKNHSelect,
	ZKNHResult
);
	input wire [63:0] A;
	input wire [3:0] ZKNHSelect;
	output wire [63:0] ZKNHResult;
	wire [31:0] sha256_32;
	wire [63:0] sha256res;
	wire [63:0] sha512res;
	sha256 sha256(
		.A(A[31:0]),
		.ZKNHSelect(ZKNHSelect[1:0]),
		.result(sha256_32)
	);
	assign sha256res = {{32 {sha256_32[31]}}, sha256_32};
	sha512_64 sha512(
		.A(A),
		.ZKNHSelect(ZKNHSelect[1:0]),
		.result(sha512res)
	);
	mux2 #(.WIDTH(64)) resultmux(
		.d0(sha256res),
		.d1(sha512res),
		.s(ZKNHSelect[3]),
		.y(ZKNHResult)
	);
endmodule
module sha256 (
	A,
	ZKNHSelect,
	result
);
	input wire [31:0] A;
	input wire [1:0] ZKNHSelect;
	output wire [31:0] result;
	wire [31:0] x [0:3][0:2];
	wire [31:0] y [0:2];
	assign x[0][0] = {A[6:0], A[31:7]};
	assign x[0][1] = {A[17:0], A[31:18]};
	assign x[0][2] = {3'b000, A[31:3]};
	assign x[1][0] = {A[16:0], A[31:17]};
	assign x[1][1] = {A[18:0], A[31:19]};
	assign x[1][2] = {10'b0000000000, A[31:10]};
	assign x[2][0] = {A[1:0], A[31:2]};
	assign x[2][1] = {A[12:0], A[31:13]};
	assign x[2][2] = {A[21:0], A[31:22]};
	assign x[3][0] = {A[5:0], A[31:6]};
	assign x[3][1] = {A[10:0], A[31:11]};
	assign x[3][2] = {A[24:0], A[31:25]};
	assign y[0] = x[ZKNHSelect[1:0]][0];
	assign y[1] = x[ZKNHSelect[1:0]][1];
	assign y[2] = x[ZKNHSelect[1:0]][2];
	assign result = (y[0] ^ y[1]) ^ y[2];
endmodule
module sha512_32 (
	A,
	B,
	ZKNHSelect,
	result
);
	input wire [31:0] A;
	input wire [31:0] B;
	input wire [2:0] ZKNHSelect;
	output wire [31:0] result;
	wire [31:0] x [0:3][0:2];
	wire [31:0] y [0:2];
	assign x[0][0] = {B[0], A[31:1]};
	assign x[0][1] = {B[7:0], A[31:8]};
	assign x[0][2] = {B[6:0] & {7 {ZKNHSelect[0]}}, A[31:7]};
	assign x[1][0] = {A[28:0], B[31:29]};
	assign x[1][1] = {B[18:0], A[31:19]};
	assign x[1][2] = {B[5:0] & {6 {ZKNHSelect[0]}}, A[31:6]};
	assign x[2][0] = {A[6:0], B[31:7]};
	assign x[2][1] = {A[1:0], B[31:2]};
	assign x[2][2] = {B[27:0], A[31:28]};
	assign x[3][0] = {A[8:0], B[31:9]};
	assign x[3][1] = {B[13:0], A[31:14]};
	assign x[3][2] = {B[17:0], A[31:18]};
	assign y[0] = x[ZKNHSelect[2:1]][0];
	assign y[1] = x[ZKNHSelect[2:1]][1];
	assign y[2] = x[ZKNHSelect[2:1]][2];
	assign result = (y[0] ^ y[1]) ^ y[2];
endmodule
module sha512_64 (
	A,
	ZKNHSelect,
	result
);
	input wire [63:0] A;
	input wire [1:0] ZKNHSelect;
	output wire [63:0] result;
	wire [63:0] x [0:3][0:2];
	wire [63:0] y [0:2];
	assign x[0][0] = {A[0], A[63:1]};
	assign x[0][1] = {A[7:0], A[63:8]};
	assign x[0][2] = {7'b0000000, A[63:7]};
	assign x[1][0] = {A[18:0], A[63:19]};
	assign x[1][1] = {A[60:0], A[63:61]};
	assign x[1][2] = {6'b000000, A[63:6]};
	assign x[2][0] = {A[27:0], A[63:28]};
	assign x[2][1] = {A[33:0], A[63:34]};
	assign x[2][2] = {A[38:0], A[63:39]};
	assign x[3][0] = {A[13:0], A[63:14]};
	assign x[3][1] = {A[17:0], A[63:18]};
	assign x[3][2] = {A[40:0], A[63:41]};
	assign y[0] = x[ZKNHSelect[1:0]][0];
	assign y[1] = x[ZKNHSelect[1:0]][1];
	assign y[2] = x[ZKNHSelect[1:0]][2];
	assign result = (y[0] ^ y[1]) ^ y[2];
endmodule
module RASPredictor (
	clk,
	reset,
	StallD,
	StallE,
	StallM,
	FlushD,
	FlushE,
	FlushM,
	BPReturnWrongD,
	ReturnD,
	ReturnE,
	CallE,
	BPReturnF,
	PCLinkE,
	RASPCF
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallD;
	input wire StallE;
	input wire StallM;
	input wire FlushD;
	input wire FlushE;
	input wire FlushM;
	input wire BPReturnWrongD;
	input wire ReturnD;
	input wire ReturnE;
	input wire CallE;
	input wire BPReturnF;
	input wire [$signed(P[4216-:32]) - 1:0] PCLinkE;
	output wire [$signed(P[4216-:32]) - 1:0] RASPCF;
	wire CounterEn;
	localparam Depth = $clog2($signed(P[1855-:32]));
	wire [Depth - 1:0] NextPtr;
	wire [Depth - 1:0] Ptr;
	wire [Depth - 1:0] P1;
	wire [Depth - 1:0] M1;
	wire [Depth - 1:0] IncDecPtr;
	reg [($signed(P[1855-:32]) * $signed(P[4216-:32])) - 1:0] memory;
	integer index;
	wire PopF;
	wire PushE;
	wire RepairD;
	wire IncrRepairD;
	wire DecRepairD;
	wire DecPtr;
	wire FlushedReturnDE;
	wire WrongPredReturnD;
	assign PopF = (BPReturnF & ~StallD) & ~FlushD;
	assign PushE = (CallE & ~StallM) & ~FlushM;
	assign WrongPredReturnD = (BPReturnWrongD & ~StallE) & ~FlushE;
	assign FlushedReturnDE = ((~StallE & FlushE) & ReturnD) | (FlushM & ReturnE);
	assign RepairD = WrongPredReturnD | FlushedReturnDE;
	assign IncrRepairD = FlushedReturnDE | (WrongPredReturnD & ~ReturnD);
	assign DecRepairD = WrongPredReturnD & ReturnD;
	assign CounterEn = (PopF | PushE) | RepairD;
	assign DecPtr = (PopF | DecRepairD) & ~IncrRepairD;
	assign P1 = 1;
	assign M1 = 1'sb1;
	mux2 #(.WIDTH(Depth)) PtrMux(
		.d0(P1),
		.d1(M1),
		.s(DecPtr),
		.y(IncDecPtr)
	);
	wire [Depth - 1:0] Sum;
	assign Sum = Ptr + IncDecPtr;
	generate
		if (|P[1823 + Depth:1824]) begin : genblk1
			assign NextPtr = (Sum >= P[1823 + Depth:1824] ? 0 : Sum);
		end
		else begin : genblk1
			assign NextPtr = Sum;
		end
	endgenerate
	flopenr #(.WIDTH(Depth)) PTR(
		.clk(clk),
		.reset(reset),
		.en(CounterEn),
		.d(NextPtr),
		.q(Ptr)
	);
	always @(posedge clk)
		if (reset)
			for (index = 0; index < $signed(P[1855-:32]); index = index + 1)
				memory[index * $signed(P[4216-:32])+:$signed(P[4216-:32])] <= {$signed(P[4216-:32]) {1'b0}};
		else if (PushE)
			memory[NextPtr * $signed(P[4216-:32])+:$signed(P[4216-:32])] <= PCLinkE;
	assign RASPCF = memory[Ptr * $signed(P[4216-:32])+:$signed(P[4216-:32])];
endmodule
module bpred (
	clk,
	reset,
	StallF,
	StallD,
	StallE,
	StallM,
	StallW,
	FlushD,
	FlushE,
	FlushM,
	FlushW,
	InstrD,
	PCNextF,
	PCPlus2or4F,
	PC1NextF,
	NextValidPCE,
	PCF,
	PCD,
	PCE,
	PCM,
	PostSpillInstrRawF,
	InstrValidD,
	InstrValidE,
	BranchD,
	BranchE,
	JumpD,
	JumpE,
	PCSrcE,
	IEUAdrE,
	IEUAdrM,
	PCLinkE,
	IClassM,
	BPWrongE,
	BPWrongM,
	BPDirWrongM,
	BTAWrongM,
	RASPredPCWrongM,
	IClassWrongM
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire StallF;
	input wire StallD;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushD;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	input wire [31:0] InstrD;
	input wire [$signed(P[4216-:32]) - 1:0] PCNextF;
	input wire [$signed(P[4216-:32]) - 1:0] PCPlus2or4F;
	output wire [$signed(P[4216-:32]) - 1:0] PC1NextF;
	output wire [$signed(P[4216-:32]) - 1:0] NextValidPCE;
	input wire [$signed(P[4216-:32]) - 1:0] PCF;
	input wire [$signed(P[4216-:32]) - 1:0] PCD;
	input wire [$signed(P[4216-:32]) - 1:0] PCE;
	input wire [$signed(P[4216-:32]) - 1:0] PCM;
	input wire [31:0] PostSpillInstrRawF;
	input wire InstrValidD;
	input wire InstrValidE;
	input wire BranchD;
	input wire BranchE;
	input wire JumpD;
	input wire JumpE;
	input wire PCSrcE;
	input wire [$signed(P[4216-:32]) - 1:0] IEUAdrE;
	input wire [$signed(P[4216-:32]) - 1:0] IEUAdrM;
	input wire [$signed(P[4216-:32]) - 1:0] PCLinkE;
	output wire [3:0] IClassM;
	output wire BPWrongE;
	output wire BPWrongM;
	output wire BPDirWrongM;
	output wire BTAWrongM;
	output wire RASPredPCWrongM;
	output wire IClassWrongM;
	wire [1:0] BPDirF;
	wire BPDirWrongE;
	wire [$signed(P[4216-:32]) - 1:0] BPBTAF;
	wire [$signed(P[4216-:32]) - 1:0] RASPCF;
	wire BPPCSrcF;
	wire [$signed(P[4216-:32]) - 1:0] BPPCF;
	wire [$signed(P[4216-:32]) - 1:0] PC0NextF;
	wire [$signed(P[4216-:32]) - 1:0] PCCorrectE;
	wire RASTargetWrongE;
	wire BTBCallF;
	wire BTBReturnF;
	wire BTBJumpF;
	wire BTBBranchF;
	wire BPBranchF;
	wire BPJumpF;
	wire BPReturnF;
	wire BPCallF;
	wire BPBranchD;
	wire BPJumpD;
	wire BPReturnD;
	wire BPCallD;
	wire ReturnD;
	wire CallD;
	wire ReturnE;
	wire CallE;
	wire BranchM;
	wire JumpM;
	wire ReturnM;
	wire CallM;
	wire BranchW;
	wire JumpW;
	wire ReturnW;
	wire CallW;
	wire BPReturnWrongD;
	wire BPBTAWrongM;
	wire PCSrcM;
	generate
		if (P[1983-:32] == 32'd0) begin : Predictor
			twoBitPredictor #(
				.P(P),
				.XLEN($signed(P[4216-:32])),
				.k($signed(P[1919-:32]))
			) DirPredictor(
				.clk(clk),
				.reset(reset),
				.StallF(StallF),
				.StallD(StallD),
				.StallE(StallE),
				.StallM(StallM),
				.StallW(StallW),
				.FlushD(FlushD),
				.FlushE(FlushE),
				.FlushM(FlushM),
				.FlushW(FlushW),
				.PCNextF(PCNextF),
				.PCM(PCM),
				.BPDirF(BPDirF),
				.BPDirWrongE(BPDirWrongE),
				.BranchE(BranchE),
				.BranchM(BranchM),
				.PCSrcE(PCSrcE)
			);
		end
		else if (P[1983-:32] == 32'd1) begin : Predictor
			gshare #(
				.P(P),
				.XLEN($signed(P[4216-:32])),
				.k($signed(P[1919-:32]))
			) DirPredictor(
				.clk(clk),
				.reset(reset),
				.StallF(StallF),
				.StallD(StallD),
				.StallE(StallE),
				.StallM(StallM),
				.StallW(StallW),
				.FlushD(FlushD),
				.FlushE(FlushE),
				.FlushM(FlushM),
				.FlushW(FlushW),
				.PCNextF(PCNextF),
				.PCF(PCF),
				.PCD(PCD),
				.PCE(PCE),
				.PCM(PCM),
				.BPDirF(BPDirF),
				.BPDirWrongE(BPDirWrongE),
				.BPBranchF(BPBranchF),
				.BranchD(BranchD),
				.BranchE(BranchE),
				.BranchM(BranchM),
				.BranchW(BranchW),
				.PCSrcE(PCSrcE)
			);
		end
		else if (P[1983-:32] == 32'd2) begin : Predictor
			gshare #(
				.P(P),
				.XLEN($signed(P[4216-:32])),
				.k($signed(P[1919-:32])),
				.TYPE(0)
			) DirPredictor(
				.clk(clk),
				.reset(reset),
				.StallF(StallF),
				.StallD(StallD),
				.StallE(StallE),
				.StallM(StallM),
				.StallW(StallW),
				.FlushD(FlushD),
				.FlushE(FlushE),
				.FlushM(FlushM),
				.FlushW(FlushW),
				.PCNextF(PCNextF),
				.PCF(PCF),
				.PCD(PCD),
				.PCE(PCE),
				.PCM(PCM),
				.BPDirF(BPDirF),
				.BPDirWrongE(BPDirWrongE),
				.BPBranchF(BPBranchF),
				.BranchD(BranchD),
				.BranchE(BranchE),
				.BranchM(BranchM),
				.BranchW(BranchW),
				.PCSrcE(PCSrcE)
			);
		end
		else if (P[1983-:32] == 32'd3) begin : Predictor
			gsharebasic #(
				.P(P),
				.XLEN($signed(P[4216-:32])),
				.k($signed(P[1919-:32]))
			) DirPredictor(
				.clk(clk),
				.reset(reset),
				.StallF(StallF),
				.StallD(StallD),
				.StallE(StallE),
				.StallM(StallM),
				.StallW(StallW),
				.FlushD(FlushD),
				.FlushE(FlushE),
				.FlushM(FlushM),
				.FlushW(FlushW),
				.PCNextF(PCNextF),
				.PCM(PCM),
				.BPDirF(BPDirF),
				.BPDirWrongE(BPDirWrongE),
				.BranchE(BranchE),
				.BranchM(BranchM),
				.PCSrcE(PCSrcE)
			);
		end
		else if (P[1983-:32] == 32'd4) begin : Predictor
			gsharebasic #(
				.P(P),
				.XLEN($signed(P[4216-:32])),
				.k($signed(P[1919-:32])),
				.TYPE(0)
			) DirPredictor(
				.clk(clk),
				.reset(reset),
				.StallF(StallF),
				.StallD(StallD),
				.StallE(StallE),
				.StallM(StallM),
				.StallW(StallW),
				.FlushD(FlushD),
				.FlushE(FlushE),
				.FlushM(FlushM),
				.FlushW(FlushW),
				.PCNextF(PCNextF),
				.PCM(PCM),
				.BPDirF(BPDirF),
				.BPDirWrongE(BPDirWrongE),
				.BranchE(BranchE),
				.BranchM(BranchM),
				.PCSrcE(PCSrcE)
			);
		end
		else if (P[1983-:32] == 32'd5) begin : Predictor
			localbpbasic #(
				.P(P),
				.XLEN($signed(P[4216-:32])),
				.m($signed(P[1951-:32])),
				.k($signed(P[1919-:32]))
			) DirPredictor(
				.clk(clk),
				.reset(reset),
				.StallF(StallF),
				.StallD(StallD),
				.StallE(StallE),
				.StallM(StallM),
				.StallW(StallW),
				.FlushD(FlushD),
				.FlushE(FlushE),
				.FlushM(FlushM),
				.FlushW(FlushW),
				.PCNextF(PCNextF),
				.PCM(PCM),
				.BPDirF(BPDirF),
				.BPDirWrongE(BPDirWrongE),
				.BranchE(BranchE),
				.BranchM(BranchM),
				.PCSrcE(PCSrcE)
			);
		end
		else if (P[1983-:32] == 32'd6) begin : Predictor
			localaheadbp #(
				.P(P),
				.XLEN($signed(P[4216-:32])),
				.m($signed(P[1951-:32])),
				.k($signed(P[1919-:32]))
			) DirPredictor(
				.clk(clk),
				.reset(reset),
				.StallF(StallF),
				.StallD(StallD),
				.StallE(StallE),
				.StallM(StallM),
				.StallW(StallW),
				.FlushD(FlushD),
				.FlushE(FlushE),
				.FlushM(FlushM),
				.FlushW(FlushW),
				.PCNextF(PCNextF),
				.PCM(PCM),
				.BPDirD(BPDirF),
				.BPDirWrongE(BPDirWrongE),
				.BranchE(BranchE),
				.BranchM(BranchM),
				.PCSrcE(PCSrcE)
			);
		end
		else if (P[1983-:32] == 32'd7) begin : Predictor
			localrepairbp #(
				.P(P),
				.XLEN($signed(P[4216-:32])),
				.m($signed(P[1951-:32])),
				.k($signed(P[1919-:32]))
			) DirPredictor(
				.clk(clk),
				.reset(reset),
				.StallF(StallF),
				.StallD(StallD),
				.StallE(StallE),
				.StallM(StallM),
				.StallW(StallW),
				.FlushD(FlushD),
				.FlushE(FlushE),
				.FlushM(FlushM),
				.FlushW(FlushW),
				.PCNextF(PCNextF),
				.PCE(PCE),
				.PCM(PCM),
				.BPDirD(BPDirF),
				.BPDirWrongE(BPDirWrongE),
				.BranchD(BranchD),
				.BranchE(BranchE),
				.BranchM(BranchM),
				.PCSrcE(PCSrcE)
			);
		end
	endgenerate
	flopenrc #(.WIDTH(1)) PCSrcMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(PCSrcE),
		.q(PCSrcM)
	);
	btb #(
		.P(P),
		.Depth($signed(P[1887-:32]))
	) TargetPredictor(
		.clk(clk),
		.reset(reset),
		.StallF(StallF),
		.StallD(StallD),
		.StallE(StallE),
		.StallM(StallM),
		.StallW(StallW),
		.FlushD(FlushD),
		.FlushE(FlushE),
		.FlushM(FlushM),
		.FlushW(FlushW),
		.PCNextF(PCNextF),
		.PCF(PCF),
		.PCD(PCD),
		.PCE(PCE),
		.PCM(PCM),
		.BPBTAF(BPBTAF),
		.BTBIClassF({BTBCallF, BTBReturnF, BTBJumpF, BTBBranchF}),
		.BPBTAWrongM(BPBTAWrongM),
		.IClassWrongM(IClassWrongM),
		.IEUAdrE(IEUAdrE),
		.IEUAdrM(IEUAdrM),
		.IClassD({CallD, ReturnD, JumpD, BranchD}),
		.IClassE({CallE, ReturnE, JumpE, BranchE}),
		.IClassM({CallM, ReturnM, JumpM, BranchM}),
		.IClassW({CallW, ReturnW, JumpW, BranchW})
	);
	icpred #(
		.P(P),
		.INSTR_CLASS_PRED(1)
	) icpred(
		.clk(clk),
		.reset(reset),
		.StallD(StallD),
		.StallE(StallE),
		.StallM(StallM),
		.StallW(StallW),
		.FlushD(FlushD),
		.FlushE(FlushE),
		.FlushM(FlushM),
		.PostSpillInstrRawF(PostSpillInstrRawF),
		.InstrD(InstrD),
		.BranchD(BranchD),
		.BranchE(BranchE),
		.JumpD(JumpD),
		.JumpE(JumpE),
		.BranchM(BranchM),
		.BranchW(BranchW),
		.JumpM(JumpM),
		.JumpW(JumpW),
		.CallD(CallD),
		.CallE(CallE),
		.CallM(CallM),
		.CallW(CallW),
		.ReturnD(ReturnD),
		.ReturnE(ReturnE),
		.ReturnM(ReturnM),
		.ReturnW(ReturnW),
		.BTBCallF(BTBCallF),
		.BTBReturnF(BTBReturnF),
		.BTBJumpF(BTBJumpF),
		.BTBBranchF(BTBBranchF),
		.BPCallF(BPCallF),
		.BPReturnF(BPReturnF),
		.BPJumpF(BPJumpF),
		.BPBranchF(BPBranchF),
		.IClassWrongM(IClassWrongM),
		.BPReturnWrongD(BPReturnWrongD)
	);
	RASPredictor #(.P(P)) RASPredictor(
		.clk(clk),
		.reset(reset),
		.StallD(StallD),
		.StallE(StallE),
		.StallM(StallM),
		.FlushD(FlushD),
		.FlushE(FlushE),
		.FlushM(FlushM),
		.BPReturnF(BPReturnF),
		.ReturnD(ReturnD),
		.ReturnE(ReturnE),
		.CallE(CallE),
		.BPReturnWrongD(BPReturnWrongD),
		.RASPCF(RASPCF),
		.PCLinkE(PCLinkE)
	);
	assign BPWrongE = ((PCCorrectE != PCD) & InstrValidE) & InstrValidD;
	flopenrc #(.WIDTH(1)) BPWrongMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(BPWrongE),
		.q(BPWrongM)
	);
	assign BPPCSrcF = (BPBranchF & BPDirF[1]) | BPJumpF;
	mux2 #(.WIDTH($signed(P[4216-:32]))) pcmuxbp(
		.d0(BPBTAF),
		.d1(RASPCF),
		.s(BPReturnF),
		.y(BPPCF)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) pcmux0(
		.d0(PCPlus2or4F),
		.d1(BPPCF),
		.s(BPPCSrcF),
		.y(PC0NextF)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) pcmux1(
		.d0(PC0NextF),
		.d1(PCCorrectE),
		.s(BPWrongE),
		.y(PC1NextF)
	);
	mux2 #(.WIDTH($signed(P[4216-:32]))) pccorrectemux(
		.d0(PCLinkE),
		.d1(IEUAdrE),
		.s(PCSrcE),
		.y(PCCorrectE)
	);
	generate
		if (1) begin : genblk2
			mux2 #(.WIDTH($signed(P[4216-:32]))) pcmuxBPWrongInvalidateFlush(
				.d0(PCE),
				.d1(PCF),
				.s(BPWrongM),
				.y(NextValidPCE)
			);
		end
		if (P[4071]) begin : genblk3
			wire [$signed(P[4216-:32]) - 1:0] RASPCD;
			wire [$signed(P[4216-:32]) - 1:0] RASPCE;
			wire RASPredPCWrongE;
			assign RASPredPCWrongE = ((RASPCE != IEUAdrE) & ReturnE) & PCSrcE;
			flopenrc #(.WIDTH($signed(P[4216-:32]))) RASTargetDReg(
				.clk(clk),
				.reset(reset),
				.clear(FlushD),
				.en(~StallD),
				.d(RASPCF),
				.q(RASPCD)
			);
			flopenrc #(.WIDTH($signed(P[4216-:32]))) RASTargetEReg(
				.clk(clk),
				.reset(reset),
				.clear(FlushE),
				.en(~StallE),
				.d(RASPCD),
				.q(RASPCE)
			);
			flopenrc #(.WIDTH(2)) BPPredWrongRegM(
				.clk(clk),
				.reset(reset),
				.clear(FlushM),
				.en(~StallM),
				.d({BPDirWrongE, RASPredPCWrongE}),
				.q({BPDirWrongM, RASPredPCWrongM})
			);
			assign BTAWrongM = BPBTAWrongM & PCSrcM;
		end
		else begin : genblk3
			assign {BTAWrongM, RASPredPCWrongM} = 0;
		end
	endgenerate
	assign IClassM = {CallM, ReturnM, JumpM, BranchM};
endmodule
module btb (
	clk,
	reset,
	StallF,
	StallD,
	StallE,
	StallM,
	StallW,
	FlushD,
	FlushE,
	FlushM,
	FlushW,
	PCNextF,
	PCF,
	PCD,
	PCE,
	PCM,
	BPBTAF,
	BTBIClassF,
	BPBTAWrongM,
	IClassWrongM,
	IEUAdrE,
	IEUAdrM,
	IClassD,
	IClassE,
	IClassM,
	IClassW
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter Depth = 10;
	input wire clk;
	input wire reset;
	input wire StallF;
	input wire StallD;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushD;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	input wire [$signed(P[4216-:32]) - 1:0] PCNextF;
	input wire [$signed(P[4216-:32]) - 1:0] PCF;
	input wire [$signed(P[4216-:32]) - 1:0] PCD;
	input wire [$signed(P[4216-:32]) - 1:0] PCE;
	input wire [$signed(P[4216-:32]) - 1:0] PCM;
	output wire [$signed(P[4216-:32]) - 1:0] BPBTAF;
	output wire [3:0] BTBIClassF;
	output wire BPBTAWrongM;
	input wire IClassWrongM;
	input wire [$signed(P[4216-:32]) - 1:0] IEUAdrE;
	input wire [$signed(P[4216-:32]) - 1:0] IEUAdrM;
	input wire [3:0] IClassD;
	input wire [3:0] IClassE;
	input wire [3:0] IClassM;
	input wire [3:0] IClassW;
	wire [Depth - 1:0] PCNextFIndex;
	wire [Depth - 1:0] PCFIndex;
	wire [Depth - 1:0] PCDIndex;
	wire [Depth - 1:0] PCEIndex;
	wire [Depth - 1:0] PCMIndex;
	wire [Depth - 1:0] PCWIndex;
	wire MatchD;
	wire MatchE;
	wire MatchM;
	wire MatchW;
	wire MatchX;
	wire [$signed(P[4216-:32]) + 3:0] ForwardBTBPredF;
	wire [$signed(P[4216-:32]) + 3:0] TableBTBPredF;
	wire [$signed(P[4216-:32]) - 1:0] IEUAdrW;
	wire [$signed(P[4216-:32]) - 1:0] PCW;
	wire [$signed(P[4216-:32]) - 1:0] BPBTAD;
	wire [$signed(P[4216-:32]) - 1:0] BPBTAE;
	wire BPBTAWrongE;
	wire BTBWrongM;
	assign PCFIndex = {PCF[Depth + 1] ^ PCF[1], PCF[Depth:2]};
	assign PCDIndex = {PCD[Depth + 1] ^ PCD[1], PCD[Depth:2]};
	assign PCEIndex = {PCE[Depth + 1] ^ PCE[1], PCE[Depth:2]};
	assign PCMIndex = {PCM[Depth + 1] ^ PCM[1], PCM[Depth:2]};
	assign PCWIndex = {PCW[Depth + 1] ^ PCW[1], PCW[Depth:2]};
	assign PCNextFIndex = {PCNextF[Depth + 1] ^ PCNextF[1], PCNextF[Depth:2]};
	assign MatchD = PCFIndex == PCDIndex;
	assign MatchE = PCFIndex == PCEIndex;
	assign MatchM = PCFIndex == PCMIndex;
	assign MatchW = PCFIndex == PCWIndex;
	assign MatchX = ((MatchD | MatchE) | MatchM) | MatchW;
	assign ForwardBTBPredF = (MatchD ? {IClassD, BPBTAD} : (MatchE ? {IClassE, IEUAdrE} : (MatchM ? {IClassM, IEUAdrM} : {IClassW, IEUAdrW})));
	assign {BTBIClassF, BPBTAF} = (MatchX ? ForwardBTBPredF : {TableBTBPredF});
	localparam sv2v_uu_memory_WIDTH = $signed(P[4216-:32]) + 4;
	localparam [(sv2v_uu_memory_WIDTH - 1) / 8:0] sv2v_uu_memory_ext_bwe2_1 = 1'sb1;
	ram2p1r1wbe #(
		.USE_SRAM(P[1743]),
		.DEPTH(2 ** Depth),
		.WIDTH($signed(P[4216-:32]) + 4)
	) memory(
		.clk(clk),
		.ce1(~StallF | reset),
		.ra1(PCNextFIndex),
		.rd1(TableBTBPredF),
		.ce2(~StallW & ~FlushW),
		.wa2(PCMIndex),
		.wd2({IClassM, IEUAdrM}),
		.we2(BTBWrongM),
		.bwe2(sv2v_uu_memory_ext_bwe2_1)
	);
	flopenrc #(.WIDTH($signed(P[4216-:32]))) BTBD(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallD),
		.d(BPBTAF),
		.q(BPBTAD)
	);
	flopenrc #(.WIDTH($signed(P[4216-:32]))) BTBTargetEReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(BPBTAD),
		.q(BPBTAE)
	);
	assign BPBTAWrongE = (BPBTAE != IEUAdrE) & (IClassE[0] | (IClassE[1] & ~IClassE[2]));
	flopenrc #(.WIDTH(1)) BPBTAWrongMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(BPBTAWrongE),
		.q(BPBTAWrongM)
	);
	assign BTBWrongM = BPBTAWrongM | IClassWrongM;
	flopenr #(.WIDTH($signed(P[4216-:32]))) PCWReg(
		.clk(clk),
		.reset(reset),
		.en(~StallW),
		.d(PCM),
		.q(PCW)
	);
	flopenr #(.WIDTH($signed(P[4216-:32]))) IEUAdrWReg(
		.clk(clk),
		.reset(reset),
		.en(~StallW),
		.d(IEUAdrM),
		.q(IEUAdrW)
	);
endmodule
module gshare (
	clk,
	reset,
	StallF,
	StallD,
	StallE,
	StallM,
	StallW,
	FlushD,
	FlushE,
	FlushM,
	FlushW,
	BPDirF,
	BPDirWrongE,
	PCNextF,
	PCF,
	PCD,
	PCE,
	PCM,
	BPBranchF,
	BranchD,
	BranchE,
	BranchM,
	BranchW,
	PCSrcE
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter XLEN = 0;
	parameter k = 10;
	parameter integer TYPE = 1;
	input wire clk;
	input wire reset;
	input wire StallF;
	input wire StallD;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushD;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	output wire [1:0] BPDirF;
	output wire BPDirWrongE;
	input wire [XLEN - 1:0] PCNextF;
	input wire [XLEN - 1:0] PCF;
	input wire [XLEN - 1:0] PCD;
	input wire [XLEN - 1:0] PCE;
	input wire [XLEN - 1:0] PCM;
	input wire BPBranchF;
	input wire BranchD;
	input wire BranchE;
	input wire BranchM;
	input wire BranchW;
	input wire PCSrcE;
	wire MatchD;
	wire MatchE;
	wire MatchM;
	wire MatchW;
	wire MatchX;
	wire [1:0] PHTBPDirF;
	wire [1:0] BPDirD;
	wire [1:0] BPDirE;
	wire [1:0] FwdNewBPDirF;
	wire [1:0] NewBPDirE;
	wire [1:0] NewBPDirM;
	wire [1:0] NewBPDirW;
	wire [k - 1:0] IndexNextF;
	wire [k - 1:0] IndexF;
	wire [k - 1:0] IndexD;
	wire [k - 1:0] IndexE;
	wire [k - 1:0] IndexM;
	wire [k - 1:0] IndexW;
	wire [k - 1:0] GHRF;
	wire [k - 1:0] GHRD;
	wire [k - 1:0] GHRE;
	wire [k - 1:0] GHRM;
	wire [k - 1:0] GHRNextM;
	wire [k - 1:0] GHRNextF;
	wire PCSrcM;
	generate
		if (TYPE == 1) begin : genblk1
			assign IndexNextF = GHRNextF ^ {PCNextF[k + 1] ^ PCNextF[1], PCNextF[k:2]};
			assign IndexF = GHRF ^ {PCF[k + 1] ^ PCF[1], PCF[k:2]};
			assign IndexD = GHRD ^ {PCD[k + 1] ^ PCD[1], PCD[k:2]};
			assign IndexE = GHRE ^ {PCE[k + 1] ^ PCE[1], PCE[k:2]};
			assign IndexM = GHRM ^ {PCM[k + 1] ^ PCM[1], PCM[k:2]};
		end
		else if (TYPE == 0) begin : genblk1
			assign IndexNextF = GHRNextF;
			assign IndexF = GHRF;
			assign IndexD = GHRD;
			assign IndexE = GHRE;
			assign IndexM = GHRM;
		end
	endgenerate
	flopenrc #(.WIDTH(k)) IndexWReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(IndexM),
		.q(IndexW)
	);
	assign MatchD = (BranchD & ~FlushE) & (IndexF == IndexD);
	assign MatchE = (BranchE & ~FlushM) & (IndexF == IndexE);
	assign MatchM = (BranchM & ~FlushW) & (IndexF == IndexM);
	assign MatchW = (BranchW & ~FlushW) & (IndexF == IndexW);
	assign MatchX = ((MatchD | MatchE) | MatchM) | MatchW;
	assign FwdNewBPDirF = (MatchD ? {2 {BPDirD[1]}} : (MatchE ? {NewBPDirE} : (MatchM ? {NewBPDirM} : NewBPDirW)));
	assign BPDirF = (MatchX ? FwdNewBPDirF : PHTBPDirF);
	ram2p1r1wbe #(
		.USE_SRAM(P[1743]),
		.DEPTH(2 ** k),
		.WIDTH(2)
	) PHT(
		.clk(clk),
		.ce1(~StallF),
		.ce2(~StallW & ~FlushW),
		.ra1(IndexNextF),
		.rd1(PHTBPDirF),
		.wa2(IndexM),
		.wd2(NewBPDirM),
		.we2(BranchM),
		.bwe2(1'b1)
	);
	flopenrc #(.WIDTH(2)) PredictionRegD(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallD),
		.d(BPDirF),
		.q(BPDirD)
	);
	flopenrc #(.WIDTH(2)) PredictionRegE(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(BPDirD),
		.q(BPDirE)
	);
	satCounter2 BPDirUpdateE(
		.BrDir(PCSrcE),
		.OldState(BPDirE),
		.NewState(NewBPDirE)
	);
	flopenrc #(.WIDTH(2)) NewPredictionRegM(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(NewBPDirE),
		.q(NewBPDirM)
	);
	flopenrc #(.WIDTH(2)) NewPredictionRegW(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(NewBPDirM),
		.q(NewBPDirW)
	);
	assign BPDirWrongE = (PCSrcE != BPDirE[1]) & BranchE;
	assign GHRNextF = (BPBranchF ? {BPDirF[1], GHRF[k - 1:1]} : GHRF);
	assign GHRF = (BranchD ? {BPDirD[1], GHRD[k - 1:1]} : GHRD);
	assign GHRD = (BranchE ? {PCSrcE, GHRE[k - 1:1]} : GHRE);
	assign GHRE = (BranchM ? {PCSrcM, GHRM[k - 1:1]} : GHRM);
	assign GHRNextM = {PCSrcM, GHRM[k - 1:1]};
	flopenr #(.WIDTH(k)) GHRReg(
		.clk(clk),
		.reset(reset),
		.en((~StallW & ~FlushW) & BranchM),
		.d(GHRNextM),
		.q(GHRM)
	);
	flopenrc #(.WIDTH(1)) PCSrcMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(PCSrcE),
		.q(PCSrcM)
	);
endmodule
module gsharebasic (
	clk,
	reset,
	StallF,
	StallD,
	StallE,
	StallM,
	StallW,
	FlushD,
	FlushE,
	FlushM,
	FlushW,
	BPDirF,
	BPDirWrongE,
	PCNextF,
	PCM,
	BranchE,
	BranchM,
	PCSrcE
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter XLEN = 0;
	parameter k = 10;
	parameter TYPE = 1;
	input wire clk;
	input wire reset;
	input wire StallF;
	input wire StallD;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushD;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	output wire [1:0] BPDirF;
	output wire BPDirWrongE;
	input wire [XLEN - 1:0] PCNextF;
	input wire [XLEN - 1:0] PCM;
	input wire BranchE;
	input wire BranchM;
	input wire PCSrcE;
	wire [k - 1:0] IndexNextF;
	wire [k - 1:0] IndexM;
	wire [1:0] BPDirD;
	wire [1:0] BPDirE;
	wire [1:0] NewBPDirE;
	wire [1:0] NewBPDirM;
	wire [k - 1:0] GHRF;
	wire [k - 1:0] GHRD;
	wire [k - 1:0] GHRE;
	wire [k - 1:0] GHRM;
	wire [k - 1:0] GHR;
	wire [k - 1:0] GHRNext;
	wire PCSrcM;
	generate
		if (TYPE == 1) begin : genblk1
			assign IndexNextF = GHR ^ {PCNextF[k + 1] ^ PCNextF[1], PCNextF[k:2]};
			assign IndexM = GHRM ^ {PCM[k + 1] ^ PCM[1], PCM[k:2]};
		end
		else if (TYPE == 0) begin : genblk1
			assign IndexNextF = GHRNext;
			assign IndexM = GHRM;
		end
	endgenerate
	ram2p1r1wbe #(
		.USE_SRAM(P[1743]),
		.DEPTH(2 ** k),
		.WIDTH(2)
	) PHT(
		.clk(clk),
		.ce1(~StallF),
		.ce2(~StallW & ~FlushW),
		.ra1(IndexNextF),
		.rd1(BPDirF),
		.wa2(IndexM),
		.wd2(NewBPDirM),
		.we2(BranchM),
		.bwe2(1'b1)
	);
	flopenrc #(.WIDTH(2)) PredictionRegD(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallD),
		.d(BPDirF),
		.q(BPDirD)
	);
	flopenrc #(.WIDTH(2)) PredictionRegE(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(BPDirD),
		.q(BPDirE)
	);
	satCounter2 BPDirUpdateE(
		.BrDir(PCSrcE),
		.OldState(BPDirE),
		.NewState(NewBPDirE)
	);
	flopenrc #(.WIDTH(2)) NewPredictionRegM(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(NewBPDirE),
		.q(NewBPDirM)
	);
	assign BPDirWrongE = (PCSrcE != BPDirE[1]) & BranchE;
	assign GHRNext = (BranchM ? {PCSrcM, GHR[k - 1:1]} : GHR);
	flopenr #(.WIDTH(k)) GHRReg(
		.clk(clk),
		.reset(reset),
		.en((~StallM & ~FlushM) & BranchM),
		.d(GHRNext),
		.q(GHR)
	);
	flopenrc #(.WIDTH(1)) PCSrcMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(PCSrcE),
		.q(PCSrcM)
	);
	flopenrc #(.WIDTH(k)) GHRFReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallF),
		.d(GHR),
		.q(GHRF)
	);
	flopenrc #(.WIDTH(k)) GHRDReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallD),
		.d(GHRF),
		.q(GHRD)
	);
	flopenrc #(.WIDTH(k)) GHREReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(GHRD),
		.q(GHRE)
	);
	flopenrc #(.WIDTH(k)) GHRMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(GHRE),
		.q(GHRM)
	);
endmodule
module icpred (
	clk,
	reset,
	StallD,
	StallE,
	StallM,
	StallW,
	FlushD,
	FlushE,
	FlushM,
	PostSpillInstrRawF,
	InstrD,
	BranchD,
	BranchE,
	JumpD,
	JumpE,
	BranchM,
	BranchW,
	JumpM,
	JumpW,
	CallD,
	CallE,
	CallM,
	CallW,
	ReturnD,
	ReturnE,
	ReturnM,
	ReturnW,
	BTBCallF,
	BTBReturnF,
	BTBJumpF,
	BTBBranchF,
	BPCallF,
	BPReturnF,
	BPJumpF,
	BPBranchF,
	IClassWrongM,
	BPReturnWrongD
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter INSTR_CLASS_PRED = 1;
	input wire clk;
	input wire reset;
	input wire StallD;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushD;
	input wire FlushE;
	input wire FlushM;
	input wire [31:0] PostSpillInstrRawF;
	input wire [31:0] InstrD;
	input wire BranchD;
	input wire BranchE;
	input wire JumpD;
	input wire JumpE;
	output wire BranchM;
	output wire BranchW;
	output wire JumpM;
	output wire JumpW;
	output wire CallD;
	output wire CallE;
	output wire CallM;
	output wire CallW;
	output wire ReturnD;
	output wire ReturnE;
	output wire ReturnM;
	output wire ReturnW;
	input wire BTBCallF;
	input wire BTBReturnF;
	input wire BTBJumpF;
	input wire BTBBranchF;
	output wire BPCallF;
	output wire BPReturnF;
	output wire BPJumpF;
	output wire BPBranchF;
	output wire IClassWrongM;
	output wire BPReturnWrongD;
	wire IClassWrongD;
	wire BPBranchD;
	wire BPJumpD;
	wire BPReturnD;
	wire BPCallD;
	wire IClassWrongE;
	generate
		if (!INSTR_CLASS_PRED) begin : DirectClassDecode
			wire cjal;
			wire cj;
			wire cjr;
			wire cjalr;
			wire CJumpF;
			wire CBranchF;
			wire NCJumpF;
			wire NCBranchF;
			if (P[1754]) begin : genblk1
				wire [4:0] CompressedOpcF;
				assign CompressedOpcF = {PostSpillInstrRawF[1:0], PostSpillInstrRawF[15:13]};
				assign cjal = (CompressedOpcF == 5'h09) & ($signed(P[4216-:32]) == 32);
				assign cj = CompressedOpcF == 5'h0d;
				assign cjr = (((CompressedOpcF == 5'h14) & ~PostSpillInstrRawF[12]) & (PostSpillInstrRawF[6:2] == 5'b00000)) & (PostSpillInstrRawF[11:7] != 5'b00000);
				assign cjalr = (((CompressedOpcF == 5'h14) & PostSpillInstrRawF[12]) & (PostSpillInstrRawF[6:2] == 5'b00000)) & (PostSpillInstrRawF[11:7] != 5'b00000);
				assign CJumpF = ((cjal | cj) | cjr) | cjalr;
				assign CBranchF = CompressedOpcF[4:1] == 4'h7;
			end
			else begin : genblk1
				assign {cjal, cj, cjr, cjalr, CJumpF, CBranchF} = 1'sb0;
			end
			assign NCJumpF = (PostSpillInstrRawF[6:0] == 7'h67) | (PostSpillInstrRawF[6:0] == 7'h6f);
			assign NCBranchF = PostSpillInstrRawF[6:0] == 7'h63;
			assign BPBranchF = NCBranchF | (P[1754] & CBranchF);
			assign BPJumpF = NCJumpF | (P[1754] & CJumpF);
			assign BPReturnF = ((NCJumpF & ((PostSpillInstrRawF[19:15] & 5'h1b) == 5'h01)) & (PostSpillInstrRawF[11:7] == 5'b00000)) | ((P[1754] & cjr) & ((PostSpillInstrRawF[11:7] & 5'h1b) == 5'h01));
			assign BPCallF = (NCJumpF & ((PostSpillInstrRawF[11:7] & 5'h1b) == 5'h01)) | (P[1754] & (cjal | (cjalr & ((PostSpillInstrRawF[11:7] & 5'h1b) == 5'h01))));
		end
		else begin : genblk1
			assign {BPCallF, BPReturnF, BPJumpF, BPBranchF} = {BTBCallF, BTBReturnF, BTBJumpF, BTBBranchF};
		end
	endgenerate
	assign ReturnD = JumpD & ((InstrD[19:15] & 5'h1b) == 5'h01);
	assign CallD = JumpD & ((InstrD[11:7] & 5'h1b) == 5'h01);
	flopenrc #(.WIDTH(2)) InstrClassRegE(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d({CallD, ReturnD}),
		.q({CallE, ReturnE})
	);
	flopenrc #(.WIDTH(4)) InstrClassRegM(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d({CallE, ReturnE, JumpE, BranchE}),
		.q({CallM, ReturnM, JumpM, BranchM})
	);
	flopenrc #(.WIDTH(4)) InstrClassRegW(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallW),
		.d({CallM, ReturnM, JumpM, BranchM}),
		.q({CallW, ReturnW, JumpW, BranchW})
	);
	flopenrc #(.WIDTH(1)) BPClassWrongRegM(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(IClassWrongE),
		.q(IClassWrongM)
	);
	flopenrc #(.WIDTH(1)) WrongInstrClassRegE(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(IClassWrongD),
		.q(IClassWrongE)
	);
	flopenrc #(.WIDTH(4)) PredInstrClassRegD(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallD),
		.d({BPCallF, BPReturnF, BPJumpF, BPBranchF}),
		.q({BPCallD, BPReturnD, BPJumpD, BPBranchD})
	);
	assign IClassWrongD = |({BPCallD, BPReturnD, BPJumpD, BPBranchD} ^ {CallD, ReturnD, JumpD, BranchD});
	assign BPReturnWrongD = BPReturnD ^ ReturnD;
endmodule
module localaheadbp (
	clk,
	reset,
	StallF,
	StallD,
	StallE,
	StallM,
	StallW,
	FlushD,
	FlushE,
	FlushM,
	FlushW,
	BPDirD,
	BPDirWrongE,
	PCNextF,
	PCM,
	BranchE,
	BranchM,
	PCSrcE
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter XLEN = 0;
	parameter m = 6;
	parameter k = 10;
	input wire clk;
	input wire reset;
	input wire StallF;
	input wire StallD;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushD;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	output wire [1:0] BPDirD;
	output wire BPDirWrongE;
	input wire [XLEN - 1:0] PCNextF;
	input wire [XLEN - 1:0] PCM;
	input wire BranchE;
	input wire BranchM;
	input wire PCSrcE;
	wire [k - 1:0] IndexNextF;
	wire [k - 1:0] IndexM;
	wire [1:0] BPDirE;
	wire [1:0] BPDirM;
	wire [1:0] NewBPDirE;
	wire [1:0] NewBPDirM;
	wire [1:0] NewBPDirW;
	wire [k - 1:0] LHRF;
	wire [k - 1:0] LHRD;
	wire [k - 1:0] LHRE;
	wire [k - 1:0] LHRM;
	wire [k - 1:0] LHRW;
	wire [k - 1:0] LHRNextF;
	wire [k - 1:0] LHRNextW;
	wire PCSrcM;
	wire [((2 ** m) * k) - 1:0] LHRArray;
	wire [m - 1:0] IndexLHRNextF;
	wire [m - 1:0] IndexLHRM;
	wire [XLEN - 1:0] PCW;
	wire UpdateM;
	assign IndexM = LHRW;
	ram2p1r1wbe #(
		.USE_SRAM(P[1743]),
		.DEPTH(2 ** k),
		.WIDTH(2)
	) PHT(
		.clk(clk),
		.ce1(~StallD),
		.ce2(~StallW & ~FlushW),
		.ra1(LHRF),
		.rd1(BPDirD),
		.wa2(IndexM),
		.wd2(NewBPDirW),
		.we2(BranchM),
		.bwe2(1'b1)
	);
	flopenrc #(.WIDTH(2)) PredictionRegE(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(BPDirD),
		.q(BPDirE)
	);
	flopenrc #(.WIDTH(2)) PredictionRegM(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(BPDirE),
		.q(BPDirM)
	);
	satCounter2 BPDirUpdateE(
		.BrDir(PCSrcE),
		.OldState(BPDirM),
		.NewState(NewBPDirM)
	);
	flopenrc #(.WIDTH(2)) NewPredictionRegW(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(NewBPDirM),
		.q(NewBPDirW)
	);
	assign BPDirWrongE = (PCSrcE != BPDirM[1]) & BranchE;
	assign LHRNextW = (BranchM ? {PCSrcM, LHRW[k - 1:1]} : LHRW);
	assign IndexLHRM = {PCW[m + 1] ^ PCW[1], PCW[m:2]};
	assign IndexLHRNextF = {PCNextF[m + 1] ^ PCNextF[1], PCNextF[m:2]};
	localparam sv2v_uu_BHT_WIDTH = k;
	localparam [(sv2v_uu_BHT_WIDTH - 1) / 8:0] sv2v_uu_BHT_ext_bwe2_1 = 1'sb1;
	ram2p1r1wbe #(
		.USE_SRAM(P[1743]),
		.DEPTH(2 ** m),
		.WIDTH(k)
	) BHT(
		.clk(clk),
		.ce1(~StallF),
		.ce2(~StallW & ~FlushW),
		.ra1(IndexLHRNextF),
		.rd1(LHRF),
		.wa2(IndexLHRM),
		.wd2(LHRNextW),
		.we2(BranchM),
		.bwe2(sv2v_uu_BHT_ext_bwe2_1)
	);
	flopenrc #(.WIDTH(1)) PCSrcMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(PCSrcE),
		.q(PCSrcM)
	);
	flopenrc #(.WIDTH(k)) LHRDReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallD),
		.d(LHRF),
		.q(LHRD)
	);
	flopenrc #(.WIDTH(k)) LHREReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(LHRD),
		.q(LHRE)
	);
	flopenrc #(.WIDTH(k)) LHRMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(LHRE),
		.q(LHRM)
	);
	flopenrc #(.WIDTH(k)) LHRWReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(LHRM),
		.q(LHRW)
	);
	flopenr #(.WIDTH(XLEN)) PCWReg(
		.clk(clk),
		.reset(reset),
		.en(~StallW),
		.d(PCM),
		.q(PCW)
	);
endmodule
module localbpbasic (
	clk,
	reset,
	StallF,
	StallD,
	StallE,
	StallM,
	StallW,
	FlushD,
	FlushE,
	FlushM,
	FlushW,
	BPDirF,
	BPDirWrongE,
	PCNextF,
	PCM,
	BranchE,
	BranchM,
	PCSrcE
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter XLEN = 0;
	parameter m = 6;
	parameter k = 10;
	input wire clk;
	input wire reset;
	input wire StallF;
	input wire StallD;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushD;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	output wire [1:0] BPDirF;
	output wire BPDirWrongE;
	input wire [XLEN - 1:0] PCNextF;
	input wire [XLEN - 1:0] PCM;
	input wire BranchE;
	input wire BranchM;
	input wire PCSrcE;
	wire [k - 1:0] IndexNextF;
	wire [k - 1:0] IndexM;
	wire [1:0] BPDirD;
	wire [1:0] BPDirE;
	wire [1:0] NewBPDirE;
	wire [1:0] NewBPDirM;
	wire [k - 1:0] LHRF;
	wire [k - 1:0] LHRD;
	wire [k - 1:0] LHRE;
	wire [k - 1:0] LHRM;
	wire [k - 1:0] LHR;
	wire [k - 1:0] LHRNextW;
	wire PCSrcM;
	wire [((2 ** m) * k) - 1:0] LHRArray;
	wire [m - 1:0] IndexLHRNextF;
	wire [m - 1:0] IndexLHRM;
	wire UpdateM;
	assign IndexNextF = LHR;
	assign IndexM = LHRM;
	ram2p1r1wbe #(
		.USE_SRAM(P[1743]),
		.DEPTH(2 ** k),
		.WIDTH(2)
	) PHT(
		.clk(clk),
		.ce1(~StallF),
		.ce2(~StallW & ~FlushW),
		.ra1(IndexNextF),
		.rd1(BPDirF),
		.wa2(IndexM),
		.wd2(NewBPDirM),
		.we2(BranchM),
		.bwe2(1'b1)
	);
	flopenrc #(.WIDTH(2)) PredictionRegD(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallD),
		.d(BPDirF),
		.q(BPDirD)
	);
	flopenrc #(.WIDTH(2)) PredictionRegE(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(BPDirD),
		.q(BPDirE)
	);
	satCounter2 BPDirUpdateE(
		.BrDir(PCSrcE),
		.OldState(BPDirE),
		.NewState(NewBPDirE)
	);
	flopenrc #(.WIDTH(2)) NewPredictionRegM(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(NewBPDirE),
		.q(NewBPDirM)
	);
	assign BPDirWrongE = (PCSrcE != BPDirE[1]) & BranchE;
	assign LHRNextW = (BranchM ? {PCSrcM, LHRM[k - 1:1]} : LHRM);
	genvar _gv_index_12;
	assign UpdateM = (BranchM & ~StallW) & ~FlushW;
	assign IndexLHRM = {PCM[m + 1] ^ PCM[1], PCM[m:2]};
	generate
		for (_gv_index_12 = 0; _gv_index_12 < (2 ** m); _gv_index_12 = _gv_index_12 + 1) begin : localhist
			localparam index = _gv_index_12;
			flopenr #(.WIDTH(k)) LocalHistoryRegister(
				.clk(clk),
				.reset(reset),
				.en(UpdateM & (index == IndexLHRM)),
				.d(LHRNextW),
				.q(LHRArray[index * k+:k])
			);
		end
	endgenerate
	assign IndexLHRNextF = {PCNextF[m + 1] ^ PCNextF[1], PCNextF[m:2]};
	assign LHR = LHRArray[IndexLHRNextF * k+:k];
	flopenrc #(.WIDTH(1)) PCSrcMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(PCSrcE),
		.q(PCSrcM)
	);
	flopenrc #(.WIDTH(k)) LHRFReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallF),
		.d(LHR),
		.q(LHRF)
	);
	flopenrc #(.WIDTH(k)) LHRDReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallD),
		.d(LHRF),
		.q(LHRD)
	);
	flopenrc #(.WIDTH(k)) LHREReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(LHRD),
		.q(LHRE)
	);
	flopenrc #(.WIDTH(k)) LHRMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(LHRE),
		.q(LHRM)
	);
endmodule
module localrepairbp (
	clk,
	reset,
	StallF,
	StallD,
	StallE,
	StallM,
	StallW,
	FlushD,
	FlushE,
	FlushM,
	FlushW,
	BPDirD,
	BPDirWrongE,
	PCNextF,
	PCE,
	PCM,
	BranchD,
	BranchE,
	BranchM,
	PCSrcE
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter XLEN = 0;
	parameter m = 6;
	parameter k = 10;
	input wire clk;
	input wire reset;
	input wire StallF;
	input wire StallD;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushD;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	output wire [1:0] BPDirD;
	output wire BPDirWrongE;
	input wire [XLEN - 1:0] PCNextF;
	input wire [XLEN - 1:0] PCE;
	input wire [XLEN - 1:0] PCM;
	input wire BranchD;
	input wire BranchE;
	input wire BranchM;
	input wire PCSrcE;
	wire [1:0] BPDirE;
	wire [1:0] BPDirM;
	wire [1:0] NewBPDirE;
	wire [1:0] NewBPDirM;
	wire [1:0] NewBPDirW;
	wire [k - 1:0] LHRF;
	wire [k - 1:0] LHRD;
	wire [k - 1:0] LHRE;
	wire [k - 1:0] LHRM;
	wire [k - 1:0] LHRW;
	wire [k - 1:0] LHRNextF;
	wire [k - 1:0] LHRNextW;
	wire PCSrcM;
	wire [((2 ** m) * k) - 1:0] LHRArray;
	wire [m - 1:0] IndexLHRNextF;
	wire [m - 1:0] IndexLHRM;
	wire [XLEN - 1:0] PCW;
	wire [k - 1:0] LHRCommittedF;
	wire [k - 1:0] LHRSpeculativeF;
	wire [m - 1:0] IndexLHRD;
	wire [k - 1:0] LHRNextE;
	reg SpeculativeFlushedF;
	ram2p1r1wbe #(
		.USE_SRAM(P[1743]),
		.DEPTH(2 ** k),
		.WIDTH(2)
	) PHT(
		.clk(clk),
		.ce1(~StallD),
		.ce2(~StallW & ~FlushW),
		.ra1(LHRF),
		.rd1(BPDirD),
		.wa2(LHRW),
		.wd2(NewBPDirW),
		.we2(BranchM),
		.bwe2(1'b1)
	);
	flopenrc #(.WIDTH(2)) PredictionRegE(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(BPDirD),
		.q(BPDirE)
	);
	flopenrc #(.WIDTH(2)) PredictionRegM(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(BPDirE),
		.q(BPDirM)
	);
	satCounter2 BPDirUpdateE(
		.BrDir(PCSrcE),
		.OldState(BPDirM),
		.NewState(NewBPDirM)
	);
	flopenrc #(.WIDTH(2)) NewPredictionRegW(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(NewBPDirM),
		.q(NewBPDirW)
	);
	assign BPDirWrongE = (PCSrcE != BPDirM[1]) & BranchE;
	assign LHRNextW = (BranchM ? {PCSrcM, LHRW[k - 1:1]} : LHRW);
	assign IndexLHRM = {PCW[m + 1] ^ PCW[1], PCW[m:2]};
	assign IndexLHRNextF = {PCNextF[m + 1] ^ PCNextF[1], PCNextF[m:2]};
	localparam sv2v_uu_BHT_WIDTH = k;
	localparam [(sv2v_uu_BHT_WIDTH - 1) / 8:0] sv2v_uu_BHT_ext_bwe2_1 = 1'sb1;
	ram2p1r1wbe #(
		.USE_SRAM(P[1743]),
		.DEPTH(2 ** m),
		.WIDTH(k)
	) BHT(
		.clk(clk),
		.ce1(~StallF),
		.ce2(~StallW & ~FlushW),
		.ra1(IndexLHRNextF),
		.rd1(LHRCommittedF),
		.wa2(IndexLHRM),
		.wd2(LHRNextW),
		.we2(BranchM),
		.bwe2(sv2v_uu_BHT_ext_bwe2_1)
	);
	assign IndexLHRD = {PCE[m + 1] ^ PCE[1], PCE[m:2]};
	assign LHRNextE = (BranchD ? {BPDirD[1], LHRE[k - 1:1]} : LHRE);
	localparam sv2v_uu_SHB_WIDTH = k;
	localparam [(sv2v_uu_SHB_WIDTH - 1) / 8:0] sv2v_uu_SHB_ext_bwe2_1 = 1'sb1;
	ram2p1r1wbe #(
		.USE_SRAM(P[1743]),
		.DEPTH(2 ** m),
		.WIDTH(k)
	) SHB(
		.clk(clk),
		.ce1(~StallF),
		.ce2(~StallE & ~FlushE),
		.ra1(IndexLHRNextF),
		.rd1(LHRSpeculativeF),
		.wa2(IndexLHRD),
		.wd2(LHRNextE),
		.we2(BranchD),
		.bwe2(sv2v_uu_SHB_ext_bwe2_1)
	);
	reg [(2 ** m) - 1:0] FlushedBits;
	always @(posedge clk) begin
		SpeculativeFlushedF <= FlushedBits[IndexLHRNextF];
		if (reset | FlushD)
			FlushedBits <= 1'sb1;
		if ((BranchD & ~StallE) & ~FlushE)
			FlushedBits[IndexLHRD] <= 1'b0;
	end
	mux2 #(.WIDTH(k)) LHRMux(
		.d0(LHRSpeculativeF),
		.d1(LHRCommittedF),
		.s(SpeculativeFlushedF),
		.y(LHRF)
	);
	flopenrc #(.WIDTH(1)) PCSrcMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(PCSrcE),
		.q(PCSrcM)
	);
	flopenrc #(.WIDTH(k)) LHRDReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallD),
		.d(LHRF),
		.q(LHRD)
	);
	flopenrc #(.WIDTH(k)) LHREReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(LHRD),
		.q(LHRE)
	);
	flopenrc #(.WIDTH(k)) LHRMReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(LHRE),
		.q(LHRM)
	);
	flopenrc #(.WIDTH(k)) LHRWReg(
		.clk(clk),
		.reset(reset),
		.clear(FlushW),
		.en(~StallW),
		.d(LHRM),
		.q(LHRW)
	);
	flopenr #(.WIDTH(XLEN)) PCWReg(
		.clk(clk),
		.reset(reset),
		.en(~StallW),
		.d(PCM),
		.q(PCW)
	);
endmodule
module satCounter2 (
	BrDir,
	OldState,
	NewState
);
	reg _sv2v_0;
	input wire BrDir;
	input wire [1:0] OldState;
	output reg [1:0] NewState;
	always @(*) begin
		if (_sv2v_0)
			;
		case (OldState)
			2'b00:
				if (BrDir)
					NewState = 2'b01;
				else
					NewState = 2'b00;
			2'b01:
				if (BrDir)
					NewState = 2'b10;
				else
					NewState = 2'b00;
			2'b10:
				if (BrDir)
					NewState = 2'b11;
				else
					NewState = 2'b01;
			2'b11:
				if (BrDir)
					NewState = 2'b11;
				else
					NewState = 2'b10;
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
module twoBitPredictor (
	clk,
	reset,
	StallF,
	StallD,
	StallE,
	StallM,
	StallW,
	FlushD,
	FlushE,
	FlushM,
	FlushW,
	PCNextF,
	PCM,
	BPDirF,
	BPDirWrongE,
	BranchE,
	BranchM,
	PCSrcE
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter XLEN = 0;
	parameter k = 10;
	input wire clk;
	input wire reset;
	input wire StallF;
	input wire StallD;
	input wire StallE;
	input wire StallM;
	input wire StallW;
	input wire FlushD;
	input wire FlushE;
	input wire FlushM;
	input wire FlushW;
	input wire [XLEN - 1:0] PCNextF;
	input wire [XLEN - 1:0] PCM;
	output wire [1:0] BPDirF;
	output wire BPDirWrongE;
	input wire BranchE;
	input wire BranchM;
	input wire PCSrcE;
	wire [k - 1:0] IndexNextF;
	wire [k - 1:0] IndexM;
	wire [1:0] PredictionMemory;
	wire DoForwarding;
	wire DoForwardingF;
	wire [1:0] BPDirD;
	wire [1:0] BPDirE;
	wire [1:0] NewBPDirE;
	wire [1:0] NewBPDirM;
	assign IndexNextF = {PCNextF[k + 1] ^ PCNextF[1], PCNextF[k:2]};
	assign IndexM = {PCM[k + 1] ^ PCM[1], PCM[k:2]};
	ram2p1r1wbe #(
		.USE_SRAM(P[1743]),
		.DEPTH(2 ** k),
		.WIDTH(2)
	) BHT(
		.clk(clk),
		.ce1(~StallF),
		.ce2(~StallW & ~FlushW),
		.ra1(IndexNextF),
		.rd1(BPDirF),
		.wa2(IndexM),
		.wd2(NewBPDirM),
		.we2(BranchM),
		.bwe2(1'b1)
	);
	flopenrc #(.WIDTH(2)) PredictionRegD(
		.clk(clk),
		.reset(reset),
		.clear(FlushD),
		.en(~StallD),
		.d(BPDirF),
		.q(BPDirD)
	);
	flopenrc #(.WIDTH(2)) PredictionRegE(
		.clk(clk),
		.reset(reset),
		.clear(FlushE),
		.en(~StallE),
		.d(BPDirD),
		.q(BPDirE)
	);
	assign BPDirWrongE = (PCSrcE != BPDirE[1]) & BranchE;
	satCounter2 BPDirUpdateE(
		.BrDir(PCSrcE),
		.OldState(BPDirE),
		.NewState(NewBPDirE)
	);
	flopenrc #(.WIDTH(2)) NewPredictionRegM(
		.clk(clk),
		.reset(reset),
		.clear(FlushM),
		.en(~StallM),
		.d(NewBPDirE),
		.q(NewBPDirM)
	);
endmodule
module tlb (
	clk,
	reset,
	SATP_MODE,
	SATP_ASID,
	STATUS_MXR,
	STATUS_SUM,
	STATUS_MPRV,
	STATUS_MPP,
	ENVCFG_PBMTE,
	ENVCFG_ADUE,
	EffectivePrivilegeModeW,
	ReadAccess,
	WriteAccess,
	CMOpM,
	DisableTranslation,
	VAdr,
	PTE,
	PageTypeWriteVal,
	TLBWrite,
	TLBFlush,
	TLBPAdr,
	TLBMiss,
	Translate,
	TLBPageFault,
	UpdateDA,
	PBMemoryType
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter TLB_ENTRIES = 8;
	parameter ITLB = 0;
	input wire clk;
	input wire reset;
	input wire [$signed(P[1608-:32]) - 1:0] SATP_MODE;
	input wire [$signed(P[1544-:32]) - 1:0] SATP_ASID;
	input wire STATUS_MXR;
	input wire STATUS_SUM;
	input wire STATUS_MPRV;
	input wire [1:0] STATUS_MPP;
	input wire ENVCFG_PBMTE;
	input wire ENVCFG_ADUE;
	input wire [1:0] EffectivePrivilegeModeW;
	input wire ReadAccess;
	input wire WriteAccess;
	input wire [3:0] CMOpM;
	input wire DisableTranslation;
	input wire [$signed(P[4216-:32]) - 1:0] VAdr;
	input wire [$signed(P[4216-:32]) - 1:0] PTE;
	input wire [1:0] PageTypeWriteVal;
	input wire TLBWrite;
	input wire TLBFlush;
	output wire [$signed(P[1640-:32]) - 1:0] TLBPAdr;
	output wire TLBMiss;
	output wire Translate;
	output wire TLBPageFault;
	output wire UpdateDA;
	output wire [1:0] PBMemoryType;
	wire [TLB_ENTRIES - 1:0] Matches;
	wire [TLB_ENTRIES - 1:0] WriteEnables;
	wire [TLB_ENTRIES - 1:0] PTE_Gs;
	wire [TLB_ENTRIES - 1:0] PTE_NAPOTs;
	wire [$signed(P[1704-:32]) - 1:0] VPN;
	wire [$signed(P[1672-:32]) - 1:0] PPN;
	wire [11:0] PTEAccessBits;
	wire [1:0] HitPageType;
	wire CAMHit;
	wire TLBHit;
	wire SV39Mode;
	wire Misaligned;
	wire MegapageMisaligned;
	wire PTE_N;
	wire NAPOT4;
	generate
		if ($signed(P[4216-:32]) == 32) begin : genblk1
			assign MegapageMisaligned = |PPN[9:0];
			assign Misaligned = (HitPageType == 2'b01) & MegapageMisaligned;
		end
		else begin : genblk1
			wire GigapageMisaligned;
			wire TerapageMisaligned;
			assign TerapageMisaligned = |PPN[26:0];
			assign GigapageMisaligned = |PPN[17:0];
			assign MegapageMisaligned = |PPN[8:0];
			assign Misaligned = (((HitPageType == 2'b11) & TerapageMisaligned) | ((HitPageType == 2'b10) & GigapageMisaligned)) | ((HitPageType == 2'b01) & MegapageMisaligned);
		end
	endgenerate
	assign VPN = VAdr[$signed(P[1704-:32]) + 11:12];
	assign NAPOT4 = PPN[3:0] == 4'b1000;
	tlbcontrol #(
		.P(P),
		.ITLB(ITLB)
	) tlbcontrol(
		.SATP_MODE(SATP_MODE),
		.VAdr(VAdr),
		.STATUS_MXR(STATUS_MXR),
		.STATUS_SUM(STATUS_SUM),
		.STATUS_MPRV(STATUS_MPRV),
		.STATUS_MPP(STATUS_MPP),
		.ENVCFG_PBMTE(ENVCFG_PBMTE),
		.ENVCFG_ADUE(ENVCFG_ADUE),
		.EffectivePrivilegeModeW(EffectivePrivilegeModeW),
		.ReadAccess(ReadAccess),
		.WriteAccess(WriteAccess),
		.CMOpM(CMOpM),
		.DisableTranslation(DisableTranslation),
		.PTEAccessBits(PTEAccessBits),
		.CAMHit(CAMHit),
		.Misaligned(Misaligned),
		.NAPOT4(NAPOT4),
		.TLBMiss(TLBMiss),
		.TLBHit(TLBHit),
		.TLBPageFault(TLBPageFault),
		.UpdateDA(UpdateDA),
		.SV39Mode(SV39Mode),
		.Translate(Translate),
		.PTE_N(PTE_N),
		.PBMemoryType(PBMemoryType)
	);
	tlblru #(.TLB_ENTRIES(TLB_ENTRIES)) lru(
		.clk(clk),
		.reset(reset),
		.TLBWrite(TLBWrite),
		.Matches(Matches),
		.TLBHit(TLBHit),
		.WriteEnables(WriteEnables)
	);
	tlbcam #(
		.P(P),
		.TLB_ENTRIES(TLB_ENTRIES),
		.KEY_BITS($signed(P[1704-:32]) + $signed(P[1544-:32])),
		.SEGMENT_BITS($signed(P[1736-:32]))
	) tlbcam(
		.clk(clk),
		.reset(reset),
		.VPN(VPN),
		.PageTypeWriteVal(PageTypeWriteVal),
		.SV39Mode(SV39Mode),
		.TLBFlush(TLBFlush),
		.WriteEnables(WriteEnables),
		.PTE_Gs(PTE_Gs),
		.PTE_NAPOTs(PTE_NAPOTs),
		.SATP_ASID(SATP_ASID),
		.Matches(Matches),
		.HitPageType(HitPageType),
		.CAMHit(CAMHit)
	);
	tlbram #(
		.P(P),
		.TLB_ENTRIES(TLB_ENTRIES)
	) tlbram(
		.clk(clk),
		.reset(reset),
		.PTE(PTE),
		.Matches(Matches),
		.WriteEnables(WriteEnables),
		.PPN(PPN),
		.PTEAccessBits(PTEAccessBits),
		.PTE_Gs(PTE_Gs),
		.PTE_NAPOTs(PTE_NAPOTs)
	);
	tlbmixer #(.P(P)) Mixer(
		.VPN(VPN),
		.PPN(PPN),
		.HitPageType(HitPageType),
		.Offset(VAdr[11:0]),
		.TLBHit(TLBHit),
		.PTE_N(PTE_N),
		.TLBPAdr(TLBPAdr)
	);
endmodule
module tlbcam (
	clk,
	reset,
	VPN,
	PageTypeWriteVal,
	SV39Mode,
	TLBFlush,
	WriteEnables,
	PTE_Gs,
	PTE_NAPOTs,
	SATP_ASID,
	Matches,
	HitPageType,
	CAMHit
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter TLB_ENTRIES = 8;
	parameter KEY_BITS = 20;
	parameter SEGMENT_BITS = 10;
	input wire clk;
	input wire reset;
	input wire [$signed(P[1704-:32]) - 1:0] VPN;
	input wire [1:0] PageTypeWriteVal;
	input wire SV39Mode;
	input wire TLBFlush;
	input wire [TLB_ENTRIES - 1:0] WriteEnables;
	input wire [TLB_ENTRIES - 1:0] PTE_Gs;
	input wire [TLB_ENTRIES - 1:0] PTE_NAPOTs;
	input wire [$signed(P[1544-:32]) - 1:0] SATP_ASID;
	output wire [TLB_ENTRIES - 1:0] Matches;
	output wire [1:0] HitPageType;
	output wire CAMHit;
	wire [(TLB_ENTRIES * 2) - 1:0] PageTypeRead;
	tlbcamline #(
		.P(P),
		.KEY_BITS(KEY_BITS),
		.SEGMENT_BITS(SEGMENT_BITS)
	) camlines[TLB_ENTRIES - 1:0](
		.clk(clk),
		.reset(reset),
		.VPN(VPN),
		.SATP_ASID(SATP_ASID),
		.SV39Mode(SV39Mode),
		.PTE_G(PTE_Gs),
		.PTE_NAPOT(PTE_NAPOTs),
		.PageTypeWriteVal(PageTypeWriteVal),
		.TLBFlush(TLBFlush),
		.WriteEnable(WriteEnables),
		.PageTypeRead(PageTypeRead),
		.Match(Matches)
	);
	assign CAMHit = |Matches & ~TLBFlush;
	or_rows #(
		.ROWS(TLB_ENTRIES),
		.COLS(2)
	) PageTypeOr(
		.a(PageTypeRead),
		.y(HitPageType)
	);
endmodule
module tlbcamline (
	clk,
	reset,
	VPN,
	SATP_ASID,
	SV39Mode,
	WriteEnable,
	PTE_G,
	PTE_NAPOT,
	PageTypeWriteVal,
	TLBFlush,
	PageTypeRead,
	Match
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter KEY_BITS = 20;
	parameter SEGMENT_BITS = 10;
	input wire clk;
	input wire reset;
	input wire [$signed(P[1704-:32]) - 1:0] VPN;
	input wire [$signed(P[1544-:32]) - 1:0] SATP_ASID;
	input wire SV39Mode;
	input wire WriteEnable;
	input wire PTE_G;
	input wire PTE_NAPOT;
	input wire [1:0] PageTypeWriteVal;
	input wire TLBFlush;
	output wire [1:0] PageTypeRead;
	output wire Match;
	wire Valid;
	wire [KEY_BITS - 1:0] Key;
	wire [1:0] PageType;
	wire [$signed(P[1544-:32]) - 1:0] Key_ASID;
	wire [SEGMENT_BITS - 1:0] Key0;
	wire [SEGMENT_BITS - 1:0] Key1;
	wire [SEGMENT_BITS - 1:0] Query0;
	wire [SEGMENT_BITS - 1:0] Query1;
	wire MatchASID;
	wire Match0;
	wire Match1;
	assign MatchASID = (SATP_ASID == Key_ASID) | PTE_G;
	generate
		if ($signed(P[4216-:32]) == 32) begin : match
			assign {Key_ASID, Key1, Key0} = Key;
			assign {Query1, Query0} = VPN;
			assign Match0 = (Query0 == Key0) | PageType[0];
			assign Match1 = Query1 == Key1;
			assign Match = ((Match0 & Match1) & MatchASID) & Valid;
		end
		else begin : match
			wire [SEGMENT_BITS - 1:0] Key2;
			wire [SEGMENT_BITS - 1:0] Key3;
			wire [SEGMENT_BITS - 1:0] Query2;
			wire [SEGMENT_BITS - 1:0] Query3;
			wire Match2;
			wire Match3;
			wire MatchNAPOT;
			assign {Query3, Query2, Query1, Query0} = VPN;
			assign {Key_ASID, Key3, Key2, Key1, Key0} = Key;
			assign MatchNAPOT = (P[4056] & PTE_NAPOT) & (Query0[SEGMENT_BITS - 1:4] == Key0[SEGMENT_BITS - 1:4]);
			assign Match0 = ((Query0 == Key0) | (PageType > 2'd0)) | MatchNAPOT;
			assign Match1 = (Query1 == Key1) | (PageType > 2'd1);
			assign Match2 = (Query2 == Key2) | (PageType > 2'd2);
			assign Match3 = (Query3 == Key3) | SV39Mode;
			assign Match = ((((Match0 & Match1) & Match2) & Match3) & MatchASID) & Valid;
		end
	endgenerate
	flopenr #(.WIDTH(2)) pagetypeflop(
		.clk(clk),
		.reset(reset),
		.en(WriteEnable),
		.d(PageTypeWriteVal),
		.q(PageType)
	);
	assign PageTypeRead = PageType & {2 {Match}};
	flopenr #(.WIDTH(1)) validbitflop(
		.clk(clk),
		.reset(reset),
		.en(WriteEnable | TLBFlush),
		.d(~TLBFlush),
		.q(Valid)
	);
	flopenr #(.WIDTH(KEY_BITS)) keyflop(
		.clk(clk),
		.reset(reset),
		.en(WriteEnable),
		.d({SATP_ASID, VPN}),
		.q(Key)
	);
endmodule
module tlbcontrol (
	SATP_MODE,
	VAdr,
	STATUS_MXR,
	STATUS_SUM,
	STATUS_MPRV,
	STATUS_MPP,
	ENVCFG_PBMTE,
	ENVCFG_ADUE,
	EffectivePrivilegeModeW,
	ReadAccess,
	WriteAccess,
	CMOpM,
	DisableTranslation,
	PTEAccessBits,
	CAMHit,
	Misaligned,
	NAPOT4,
	TLBMiss,
	TLBHit,
	TLBPageFault,
	UpdateDA,
	SV39Mode,
	Translate,
	PTE_N,
	PBMemoryType
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter [4216:0] ITLB = 0;
	input wire [$signed(P[1608-:32]) - 1:0] SATP_MODE;
	input wire [$signed(P[4216-:32]) - 1:0] VAdr;
	input wire STATUS_MXR;
	input wire STATUS_SUM;
	input wire STATUS_MPRV;
	input wire [1:0] STATUS_MPP;
	input wire ENVCFG_PBMTE;
	input wire ENVCFG_ADUE;
	input wire [1:0] EffectivePrivilegeModeW;
	input wire ReadAccess;
	input wire WriteAccess;
	input wire [3:0] CMOpM;
	input wire DisableTranslation;
	input wire [11:0] PTEAccessBits;
	input wire CAMHit;
	input wire Misaligned;
	input wire NAPOT4;
	output wire TLBMiss;
	output wire TLBHit;
	output wire TLBPageFault;
	output wire UpdateDA;
	output wire SV39Mode;
	output wire Translate;
	output wire PTE_N;
	output wire [1:0] PBMemoryType;
	wire [1:0] PTE_PBMT;
	wire PTE_RESERVED;
	wire PTE_D;
	wire PTE_A;
	wire PTE_U;
	wire PTE_X;
	wire PTE_W;
	wire PTE_R;
	wire PTE_V;
	wire UpperBitsUnequal;
	wire TLBAccess;
	wire ImproperPrivilege;
	wire BadPBMT;
	wire BadNAPOT;
	wire BadReserved;
	wire ReservedRW;
	wire InvalidAccess;
	wire PreUpdateDA;
	wire PrePageFault;
	assign Translate = ((SATP_MODE != P[1508 + $signed(P[1608-:32]):1509]) & (EffectivePrivilegeModeW != P[1742-:2])) & ~DisableTranslation;
	assign TLBAccess = (ReadAccess | WriteAccess) | (|CMOpM);
	vm64check #(.P(P)) vm64check(
		.SATP_MODE(SATP_MODE),
		.VAdr(VAdr),
		.SV39Mode(SV39Mode),
		.UpperBitsUnequal(UpperBitsUnequal)
	);
	assign PTE_N = PTEAccessBits[11];
	assign PTE_PBMT = PTEAccessBits[10:9];
	assign PTE_RESERVED = PTEAccessBits[8];
	assign {PTE_D, PTE_A} = PTEAccessBits[7:6];
	assign {PTE_U, PTE_X, PTE_W, PTE_R, PTE_V} = PTEAccessBits[4:0];
	assign PBMemoryType = PTE_PBMT & {2 {(Translate & TLBHit) & P[4057]}};
	assign BadPBMT = ((PTE_PBMT != 0) & ~(P[4057] & ENVCFG_PBMTE)) | (PTE_PBMT == 3);
	assign BadNAPOT = PTE_N & (~P[4056] | ~NAPOT4);
	assign BadReserved = PTE_RESERVED;
	assign ReservedRW = PTE_W & ~PTE_R;
	generate
		if (ITLB == 1) begin : itlb
			assign ImproperPrivilege = ((EffectivePrivilegeModeW == P[1738-:2]) & ~PTE_U) | ((EffectivePrivilegeModeW == P[1740-:2]) & PTE_U);
			assign PreUpdateDA = ~PTE_A;
			assign InvalidAccess = ~PTE_X | ReservedRW;
		end
		else begin : dtlb
			wire InvalidRead;
			wire InvalidWrite;
			wire InvalidCBOM;
			wire InvalidCBOZ;
			assign ImproperPrivilege = ((EffectivePrivilegeModeW == P[1738-:2]) & ~PTE_U) | (((EffectivePrivilegeModeW == P[1740-:2]) & PTE_U) & ~STATUS_SUM);
			assign InvalidRead = (ReadAccess & ~PTE_R) & (~STATUS_MXR | ~PTE_X);
			assign InvalidWrite = WriteAccess & ~PTE_W;
			assign InvalidCBOM = |CMOpM[2:0] & (~PTE_R & (~STATUS_MXR | ~PTE_X));
			assign InvalidCBOZ = CMOpM[3] & ~PTE_W;
			assign InvalidAccess = (((InvalidRead | InvalidWrite) | InvalidCBOM) | InvalidCBOZ) | ReservedRW;
			assign PreUpdateDA = ~PTE_A | (WriteAccess & ~PTE_D);
		end
	endgenerate
	assign UpdateDA = ((((P[4064] & PreUpdateDA) & Translate) & TLBHit) & ~TLBPageFault) & ENVCFG_ADUE;
	assign PrePageFault = ((((UpperBitsUnequal | Misaligned) | ~PTE_V) | ImproperPrivilege) | (($signed(P[4216-:32]) == 64) & ((BadPBMT | BadNAPOT) | BadReserved))) | (PreUpdateDA & (~P[4064] | ~ENVCFG_ADUE));
	assign TLBPageFault = (Translate & TLBHit) & (PrePageFault | InvalidAccess);
	assign TLBHit = CAMHit & TLBAccess;
	assign TLBMiss = (~CAMHit & TLBAccess) & Translate;
endmodule
module tlblru (
	clk,
	reset,
	TLBWrite,
	Matches,
	TLBHit,
	WriteEnables
);
	parameter TLB_ENTRIES = 8;
	input wire clk;
	input wire reset;
	input wire TLBWrite;
	input wire [TLB_ENTRIES - 1:0] Matches;
	input wire TLBHit;
	output wire [TLB_ENTRIES - 1:0] WriteEnables;
	wire [TLB_ENTRIES - 1:0] RUBits;
	wire [TLB_ENTRIES - 1:0] RUBitsNext;
	wire [TLB_ENTRIES - 1:0] RUBitsAccessed;
	wire [TLB_ENTRIES - 1:0] WriteLines;
	wire [TLB_ENTRIES - 1:0] AccessLines;
	wire AllUsed;
	priorityonehot #(.N(TLB_ENTRIES)) nru(
		.a(~RUBits),
		.y(WriteLines)
	);
	assign WriteEnables = WriteLines & {TLB_ENTRIES {TLBWrite}};
	assign AccessLines = (TLBWrite ? WriteLines : Matches);
	assign RUBitsAccessed = AccessLines | RUBits;
	assign AllUsed = &RUBitsAccessed;
	assign RUBitsNext = (AllUsed ? 0 : RUBitsAccessed);
	flopenr #(.WIDTH(TLB_ENTRIES)) lrustate(
		.clk(clk),
		.reset(reset),
		.en(TLBHit | TLBWrite),
		.d(RUBitsNext),
		.q(RUBits)
	);
endmodule
module tlbmixer (
	VPN,
	PPN,
	HitPageType,
	Offset,
	TLBHit,
	PTE_N,
	TLBPAdr
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[1704-:32]) - 1:0] VPN;
	input wire [$signed(P[1672-:32]) - 1:0] PPN;
	input wire [1:0] HitPageType;
	input wire [11:0] Offset;
	input wire TLBHit;
	input wire PTE_N;
	output wire [$signed(P[1640-:32]) - 1:0] TLBPAdr;
	localparam EXTRA_BITS = $signed(P[1672-:32]) - $signed(P[1704-:32]);
	wire [$signed(P[1672-:32]) - 1:0] ZeroExtendedVPN;
	wire [$signed(P[1672-:32]) - 1:0] PageNumberMask;
	wire [$signed(P[1672-:32]) - 1:0] PPNMixed;
	wire [$signed(P[1672-:32]) - 1:0] PPNMixed2;
	generate
		if ($signed(P[4216-:32]) == 32) begin : genblk1
			mux2 #(.WIDTH(22)) pnm(
				.d0(22'h000000),
				.d1(22'h0003ff),
				.s(HitPageType[0]),
				.y(PageNumberMask)
			);
		end
		else begin : genblk1
			mux4 #(.WIDTH(44)) pnm(
				.d0(44'h00000000000),
				.d1(44'h000000001ff),
				.d2(44'h0000003ffff),
				.d3(44'h00007ffffff),
				.s(HitPageType),
				.y(PageNumberMask)
			);
		end
	endgenerate
	assign ZeroExtendedVPN = {{EXTRA_BITS {1'b0}}, VPN};
	assign PPNMixed = PPN | (ZeroExtendedVPN & PageNumberMask);
	generate
		if (P[4056]) begin : genblk2
			wire [3:0] PPNMixedBot;
			mux2 #(.WIDTH(4)) napotmux(
				.d0(PPNMixed[3:0]),
				.d1(VPN[3:0]),
				.s(PTE_N),
				.y(PPNMixedBot)
			);
			assign PPNMixed2 = {PPNMixed[$signed(P[1672-:32]) - 1:4], PPNMixedBot};
		end
		else begin : genblk2
			assign PPNMixed2 = PPNMixed;
		end
	endgenerate
	assign TLBPAdr = (TLBHit ? {PPNMixed2, Offset} : 0);
endmodule
module tlbram (
	clk,
	reset,
	PTE,
	Matches,
	WriteEnables,
	PPN,
	PTEAccessBits,
	PTE_Gs,
	PTE_NAPOTs
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	parameter TLB_ENTRIES = 8;
	input wire clk;
	input wire reset;
	input wire [$signed(P[4216-:32]) - 1:0] PTE;
	input wire [TLB_ENTRIES - 1:0] Matches;
	input wire [TLB_ENTRIES - 1:0] WriteEnables;
	output wire [$signed(P[1672-:32]) - 1:0] PPN;
	output wire [11:0] PTEAccessBits;
	output wire [TLB_ENTRIES - 1:0] PTE_Gs;
	output wire [TLB_ENTRIES - 1:0] PTE_NAPOTs;
	wire [(TLB_ENTRIES * $signed(P[4216-:32])) - 1:0] RamRead;
	wire [$signed(P[4216-:32]) - 1:0] PageTableEntry;
	tlbramline #(.P(P)) tlbramline[TLB_ENTRIES - 1:0](
		.clk(clk),
		.reset(reset),
		.re(Matches),
		.we(WriteEnables),
		.d(PTE),
		.q(RamRead),
		.PTE_G(PTE_Gs),
		.PTE_NAPOT(PTE_NAPOTs)
	);
	or_rows #(
		.ROWS(TLB_ENTRIES),
		.COLS($signed(P[4216-:32]))
	) PTEOr(
		.a(RamRead),
		.y(PageTableEntry)
	);
	assign PTEAccessBits = {PageTableEntry[$signed(P[4216-:32]) - 1:$signed(P[4216-:32]) - 4] & {4 {$signed(P[4216-:32]) == 64}}, PageTableEntry[7:0]};
	assign PPN = PageTableEntry[$signed(P[1672-:32]) + 9:10];
endmodule
module tlbramline (
	clk,
	reset,
	re,
	we,
	d,
	q,
	PTE_G,
	PTE_NAPOT
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire clk;
	input wire reset;
	input wire re;
	input wire we;
	input wire [$signed(P[4216-:32]) - 1:0] d;
	output wire [$signed(P[4216-:32]) - 1:0] q;
	output wire PTE_G;
	output wire PTE_NAPOT;
	wire [$signed(P[4216-:32]) - 1:0] line;
	generate
		if ($signed(P[4216-:32]) == 64) begin : genblk1
			wire [57:0] ptereg;
			wire reserved;
			assign reserved = |d[60:54];
			flopenr #(.WIDTH(58)) pteflop(
				.clk(clk),
				.reset(reset),
				.en(we),
				.d({d[63:61], reserved, d[53:0]}),
				.q(ptereg)
			);
			assign line = {ptereg[57:54], 6'b000000, ptereg[53:0]};
		end
		else begin : genblk1
			flopenr #(.WIDTH($signed(P[4216-:32]))) pteflop(
				.clk(clk),
				.reset(reset),
				.en(we),
				.d(d),
				.q(line)
			);
		end
	endgenerate
	assign q = (re ? line : 0);
	assign PTE_G = line[5];
	assign PTE_NAPOT = (P[4056] & line[$signed(P[4216-:32]) - 1]) & (line[13:10] == 4'b1000);
endmodule
module vm64check (
	SATP_MODE,
	VAdr,
	SV39Mode,
	UpperBitsUnequal
);
	parameter [4216:0] P = 4217'b00000000000000000000000001000000000000000000101000001000100101111000000000000000000000000010000000000000000000000000000000000000011100000010000011111111111111111111111000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111110100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000010000000000000000000000000000101010000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000100110000000000000000000000000000000100000000000000000000000000000110000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000001001111111011111110110100000000000000000000000000000010010000000000000000000000000010010000000000000000000000000000101100000000000000000000000000001110000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000100000000000110001001111101110110000000000000000000000000000011000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000111100000000000000000000000001110000000000000000000000111111111111111100000000000000000000000001000000000000000000000000000000000010110000000000000000000000000011010000000000000000000000001111111111010000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000111111100000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010000000000000000000000000000011111000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000101100000000000000000000000000110100010000000000000000000000111111111100000000000000000000000000000011000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000101110000000000000000000000000001111111000000000000000000000000000100000000000000000000000000000000010100000000000000000000000000001010100000000000000000000000000000111100000000000000000000000001010100000000000000000000000000010000000000000000000000000000000000011100000000000000000000000010100100000000000000000000000000000010000000000000000000000000001010001000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000100100000000000000000000000000000100000000000000000000000000010001100000000000000000000000000000011100000000000000000000000001000110;
	input wire [$signed(P[1608-:32]) - 1:0] SATP_MODE;
	input wire [$signed(P[4216-:32]) - 1:0] VAdr;
	output wire SV39Mode;
	output wire UpperBitsUnequal;
	generate
		if ($signed(P[4216-:32]) == 64) begin : genblk1
			assign SV39Mode = SATP_MODE == P[1504-:4];
			wire eq_63_47;
			wire eq_46_38;
			assign eq_46_38 = &VAdr[46:38] | ~|VAdr[46:38];
			assign eq_63_47 = &VAdr[63:47] | ~|VAdr[63:47];
			assign UpperBitsUnequal = (SV39Mode ? ~(eq_63_47 & eq_46_38) : ~eq_63_47);
		end
		else begin : genblk1
			assign SV39Mode = 1'b0;
			assign UpperBitsUnequal = 1'b0;
		end
	endgenerate
endmodule
